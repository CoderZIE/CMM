// Verilog module
module matrix_mult_optimized_10x64_8_1449#(
    parameter ROWS = 10,
    parameter COLS = 64,
    parameter MEM_SIZE = 1449,
    parameter input_bit_width = 9,
    parameter output_bit_width = 22
)(
    input wire signed [input_bit_width-1:0] input_vector [0: COLS-1],
   output wire signed [output_bit_width-1:0] output_vector [0: ROWS-1]
);

wire signed [output_bit_width-1:0] MEM [0:MEM_SIZE];

assign MEM[0] = -(input_vector[0] << 7);
assign MEM[1] = input_vector[0] << 6;
assign MEM[2] = input_vector[0] << 5;
assign MEM[3] = input_vector[0] << 4;
assign MEM[4] = input_vector[0] << 3;
assign MEM[5] = input_vector[0] << 2;
assign MEM[6] = input_vector[0] << 1;
assign MEM[7] = input_vector[0] << 0;
assign MEM[8] = -(input_vector[1] << 7);
assign MEM[9] = input_vector[1] << 6;
assign MEM[10] = input_vector[1] << 5;
assign MEM[11] = input_vector[1] << 4;
assign MEM[12] = input_vector[1] << 3;
assign MEM[13] = input_vector[1] << 2;
assign MEM[14] = input_vector[1] << 1;
assign MEM[15] = input_vector[1] << 0;
assign MEM[16] = -(input_vector[2] << 7);
assign MEM[17] = input_vector[2] << 6;
assign MEM[18] = input_vector[2] << 5;
assign MEM[19] = input_vector[2] << 4;
assign MEM[20] = input_vector[2] << 3;
assign MEM[21] = input_vector[2] << 2;
assign MEM[22] = input_vector[2] << 1;
assign MEM[23] = input_vector[2] << 0;
assign MEM[24] = -(input_vector[3] << 7);
assign MEM[25] = input_vector[3] << 6;
assign MEM[26] = input_vector[3] << 5;
assign MEM[27] = input_vector[3] << 4;
assign MEM[28] = input_vector[3] << 3;
assign MEM[29] = input_vector[3] << 2;
assign MEM[30] = input_vector[3] << 1;
assign MEM[31] = input_vector[3] << 0;
assign MEM[32] = -(input_vector[4] << 7);
assign MEM[33] = input_vector[4] << 6;
assign MEM[34] = input_vector[4] << 5;
assign MEM[35] = input_vector[4] << 4;
assign MEM[36] = input_vector[4] << 3;
assign MEM[37] = input_vector[4] << 2;
assign MEM[38] = input_vector[4] << 1;
assign MEM[39] = input_vector[4] << 0;
assign MEM[40] = -(input_vector[5] << 7);
assign MEM[41] = input_vector[5] << 6;
assign MEM[42] = input_vector[5] << 5;
assign MEM[43] = input_vector[5] << 4;
assign MEM[44] = input_vector[5] << 3;
assign MEM[45] = input_vector[5] << 2;
assign MEM[46] = input_vector[5] << 1;
assign MEM[47] = input_vector[5] << 0;
assign MEM[48] = -(input_vector[6] << 7);
assign MEM[49] = input_vector[6] << 6;
assign MEM[50] = input_vector[6] << 5;
assign MEM[51] = input_vector[6] << 4;
assign MEM[52] = input_vector[6] << 3;
assign MEM[53] = input_vector[6] << 2;
assign MEM[54] = input_vector[6] << 1;
assign MEM[55] = input_vector[6] << 0;
assign MEM[56] = -(input_vector[7] << 7);
assign MEM[57] = input_vector[7] << 6;
assign MEM[58] = input_vector[7] << 5;
assign MEM[59] = input_vector[7] << 4;
assign MEM[60] = input_vector[7] << 3;
assign MEM[61] = input_vector[7] << 2;
assign MEM[62] = input_vector[7] << 1;
assign MEM[63] = input_vector[7] << 0;
assign MEM[64] = -(input_vector[8] << 7);
assign MEM[65] = input_vector[8] << 6;
assign MEM[66] = input_vector[8] << 5;
assign MEM[67] = input_vector[8] << 4;
assign MEM[68] = input_vector[8] << 3;
assign MEM[69] = input_vector[8] << 2;
assign MEM[70] = input_vector[8] << 1;
assign MEM[71] = input_vector[8] << 0;
assign MEM[72] = -(input_vector[9] << 7);
assign MEM[73] = input_vector[9] << 6;
assign MEM[74] = input_vector[9] << 5;
assign MEM[75] = input_vector[9] << 4;
assign MEM[76] = input_vector[9] << 3;
assign MEM[77] = input_vector[9] << 2;
assign MEM[78] = input_vector[9] << 1;
assign MEM[79] = input_vector[9] << 0;
assign MEM[80] = -(input_vector[10] << 7);
assign MEM[81] = input_vector[10] << 6;
assign MEM[82] = input_vector[10] << 5;
assign MEM[83] = input_vector[10] << 4;
assign MEM[84] = input_vector[10] << 3;
assign MEM[85] = input_vector[10] << 2;
assign MEM[86] = input_vector[10] << 1;
assign MEM[87] = input_vector[10] << 0;
assign MEM[88] = -(input_vector[11] << 7);
assign MEM[89] = input_vector[11] << 6;
assign MEM[90] = input_vector[11] << 5;
assign MEM[91] = input_vector[11] << 4;
assign MEM[92] = input_vector[11] << 3;
assign MEM[93] = input_vector[11] << 2;
assign MEM[94] = input_vector[11] << 1;
assign MEM[95] = input_vector[11] << 0;
assign MEM[96] = -(input_vector[12] << 7);
assign MEM[97] = input_vector[12] << 6;
assign MEM[98] = input_vector[12] << 5;
assign MEM[99] = input_vector[12] << 4;
assign MEM[100] = input_vector[12] << 3;
assign MEM[101] = input_vector[12] << 2;
assign MEM[102] = input_vector[12] << 1;
assign MEM[103] = input_vector[12] << 0;
assign MEM[104] = -(input_vector[13] << 7);
assign MEM[105] = input_vector[13] << 6;
assign MEM[106] = input_vector[13] << 5;
assign MEM[107] = input_vector[13] << 4;
assign MEM[108] = input_vector[13] << 3;
assign MEM[109] = input_vector[13] << 2;
assign MEM[110] = input_vector[13] << 1;
assign MEM[111] = input_vector[13] << 0;
assign MEM[112] = -(input_vector[14] << 7);
assign MEM[113] = input_vector[14] << 6;
assign MEM[114] = input_vector[14] << 5;
assign MEM[115] = input_vector[14] << 4;
assign MEM[116] = input_vector[14] << 3;
assign MEM[117] = input_vector[14] << 2;
assign MEM[118] = input_vector[14] << 1;
assign MEM[119] = input_vector[14] << 0;
assign MEM[120] = -(input_vector[15] << 7);
assign MEM[121] = input_vector[15] << 6;
assign MEM[122] = input_vector[15] << 5;
assign MEM[123] = input_vector[15] << 4;
assign MEM[124] = input_vector[15] << 3;
assign MEM[125] = input_vector[15] << 2;
assign MEM[126] = input_vector[15] << 1;
assign MEM[127] = input_vector[15] << 0;
assign MEM[128] = -(input_vector[16] << 7);
assign MEM[129] = input_vector[16] << 6;
assign MEM[130] = input_vector[16] << 5;
assign MEM[131] = input_vector[16] << 4;
assign MEM[132] = input_vector[16] << 3;
assign MEM[133] = input_vector[16] << 2;
assign MEM[134] = input_vector[16] << 1;
assign MEM[135] = input_vector[16] << 0;
assign MEM[136] = -(input_vector[17] << 7);
assign MEM[137] = input_vector[17] << 6;
assign MEM[138] = input_vector[17] << 5;
assign MEM[139] = input_vector[17] << 4;
assign MEM[140] = input_vector[17] << 3;
assign MEM[141] = input_vector[17] << 2;
assign MEM[142] = input_vector[17] << 1;
assign MEM[143] = input_vector[17] << 0;
assign MEM[144] = -(input_vector[18] << 7);
assign MEM[145] = input_vector[18] << 6;
assign MEM[146] = input_vector[18] << 5;
assign MEM[147] = input_vector[18] << 4;
assign MEM[148] = input_vector[18] << 3;
assign MEM[149] = input_vector[18] << 2;
assign MEM[150] = input_vector[18] << 1;
assign MEM[151] = input_vector[18] << 0;
assign MEM[152] = -(input_vector[19] << 7);
assign MEM[153] = input_vector[19] << 6;
assign MEM[154] = input_vector[19] << 5;
assign MEM[155] = input_vector[19] << 4;
assign MEM[156] = input_vector[19] << 3;
assign MEM[157] = input_vector[19] << 2;
assign MEM[158] = input_vector[19] << 1;
assign MEM[159] = input_vector[19] << 0;
assign MEM[160] = -(input_vector[20] << 7);
assign MEM[161] = input_vector[20] << 6;
assign MEM[162] = input_vector[20] << 5;
assign MEM[163] = input_vector[20] << 4;
assign MEM[164] = input_vector[20] << 3;
assign MEM[165] = input_vector[20] << 2;
assign MEM[166] = input_vector[20] << 1;
assign MEM[167] = input_vector[20] << 0;
assign MEM[168] = -(input_vector[21] << 7);
assign MEM[169] = input_vector[21] << 6;
assign MEM[170] = input_vector[21] << 5;
assign MEM[171] = input_vector[21] << 4;
assign MEM[172] = input_vector[21] << 3;
assign MEM[173] = input_vector[21] << 2;
assign MEM[174] = input_vector[21] << 1;
assign MEM[175] = input_vector[21] << 0;
assign MEM[176] = -(input_vector[22] << 7);
assign MEM[177] = input_vector[22] << 6;
assign MEM[178] = input_vector[22] << 5;
assign MEM[179] = input_vector[22] << 4;
assign MEM[180] = input_vector[22] << 3;
assign MEM[181] = input_vector[22] << 2;
assign MEM[182] = input_vector[22] << 1;
assign MEM[183] = input_vector[22] << 0;
assign MEM[184] = -(input_vector[23] << 7);
assign MEM[185] = input_vector[23] << 6;
assign MEM[186] = input_vector[23] << 5;
assign MEM[187] = input_vector[23] << 4;
assign MEM[188] = input_vector[23] << 3;
assign MEM[189] = input_vector[23] << 2;
assign MEM[190] = input_vector[23] << 1;
assign MEM[191] = input_vector[23] << 0;
assign MEM[192] = -(input_vector[24] << 7);
assign MEM[193] = input_vector[24] << 6;
assign MEM[194] = input_vector[24] << 5;
assign MEM[195] = input_vector[24] << 4;
assign MEM[196] = input_vector[24] << 3;
assign MEM[197] = input_vector[24] << 2;
assign MEM[198] = input_vector[24] << 1;
assign MEM[199] = input_vector[24] << 0;
assign MEM[200] = -(input_vector[25] << 7);
assign MEM[201] = input_vector[25] << 6;
assign MEM[202] = input_vector[25] << 5;
assign MEM[203] = input_vector[25] << 4;
assign MEM[204] = input_vector[25] << 3;
assign MEM[205] = input_vector[25] << 2;
assign MEM[206] = input_vector[25] << 1;
assign MEM[207] = input_vector[25] << 0;
assign MEM[208] = -(input_vector[26] << 7);
assign MEM[209] = input_vector[26] << 6;
assign MEM[210] = input_vector[26] << 5;
assign MEM[211] = input_vector[26] << 4;
assign MEM[212] = input_vector[26] << 3;
assign MEM[213] = input_vector[26] << 2;
assign MEM[214] = input_vector[26] << 1;
assign MEM[215] = input_vector[26] << 0;
assign MEM[216] = -(input_vector[27] << 7);
assign MEM[217] = input_vector[27] << 6;
assign MEM[218] = input_vector[27] << 5;
assign MEM[219] = input_vector[27] << 4;
assign MEM[220] = input_vector[27] << 3;
assign MEM[221] = input_vector[27] << 2;
assign MEM[222] = input_vector[27] << 1;
assign MEM[223] = input_vector[27] << 0;
assign MEM[224] = -(input_vector[28] << 7);
assign MEM[225] = input_vector[28] << 6;
assign MEM[226] = input_vector[28] << 5;
assign MEM[227] = input_vector[28] << 4;
assign MEM[228] = input_vector[28] << 3;
assign MEM[229] = input_vector[28] << 2;
assign MEM[230] = input_vector[28] << 1;
assign MEM[231] = input_vector[28] << 0;
assign MEM[232] = -(input_vector[29] << 7);
assign MEM[233] = input_vector[29] << 6;
assign MEM[234] = input_vector[29] << 5;
assign MEM[235] = input_vector[29] << 4;
assign MEM[236] = input_vector[29] << 3;
assign MEM[237] = input_vector[29] << 2;
assign MEM[238] = input_vector[29] << 1;
assign MEM[239] = input_vector[29] << 0;
assign MEM[240] = -(input_vector[30] << 7);
assign MEM[241] = input_vector[30] << 6;
assign MEM[242] = input_vector[30] << 5;
assign MEM[243] = input_vector[30] << 4;
assign MEM[244] = input_vector[30] << 3;
assign MEM[245] = input_vector[30] << 2;
assign MEM[246] = input_vector[30] << 1;
assign MEM[247] = input_vector[30] << 0;
assign MEM[248] = -(input_vector[31] << 7);
assign MEM[249] = input_vector[31] << 6;
assign MEM[250] = input_vector[31] << 5;
assign MEM[251] = input_vector[31] << 4;
assign MEM[252] = input_vector[31] << 3;
assign MEM[253] = input_vector[31] << 2;
assign MEM[254] = input_vector[31] << 1;
assign MEM[255] = input_vector[31] << 0;
assign MEM[256] = -(input_vector[32] << 7);
assign MEM[257] = input_vector[32] << 6;
assign MEM[258] = input_vector[32] << 5;
assign MEM[259] = input_vector[32] << 4;
assign MEM[260] = input_vector[32] << 3;
assign MEM[261] = input_vector[32] << 2;
assign MEM[262] = input_vector[32] << 1;
assign MEM[263] = input_vector[32] << 0;
assign MEM[264] = -(input_vector[33] << 7);
assign MEM[265] = input_vector[33] << 6;
assign MEM[266] = input_vector[33] << 5;
assign MEM[267] = input_vector[33] << 4;
assign MEM[268] = input_vector[33] << 3;
assign MEM[269] = input_vector[33] << 2;
assign MEM[270] = input_vector[33] << 1;
assign MEM[271] = input_vector[33] << 0;
assign MEM[272] = -(input_vector[34] << 7);
assign MEM[273] = input_vector[34] << 6;
assign MEM[274] = input_vector[34] << 5;
assign MEM[275] = input_vector[34] << 4;
assign MEM[276] = input_vector[34] << 3;
assign MEM[277] = input_vector[34] << 2;
assign MEM[278] = input_vector[34] << 1;
assign MEM[279] = input_vector[34] << 0;
assign MEM[280] = -(input_vector[35] << 7);
assign MEM[281] = input_vector[35] << 6;
assign MEM[282] = input_vector[35] << 5;
assign MEM[283] = input_vector[35] << 4;
assign MEM[284] = input_vector[35] << 3;
assign MEM[285] = input_vector[35] << 2;
assign MEM[286] = input_vector[35] << 1;
assign MEM[287] = input_vector[35] << 0;
assign MEM[288] = -(input_vector[36] << 7);
assign MEM[289] = input_vector[36] << 6;
assign MEM[290] = input_vector[36] << 5;
assign MEM[291] = input_vector[36] << 4;
assign MEM[292] = input_vector[36] << 3;
assign MEM[293] = input_vector[36] << 2;
assign MEM[294] = input_vector[36] << 1;
assign MEM[295] = input_vector[36] << 0;
assign MEM[296] = -(input_vector[37] << 7);
assign MEM[297] = input_vector[37] << 6;
assign MEM[298] = input_vector[37] << 5;
assign MEM[299] = input_vector[37] << 4;
assign MEM[300] = input_vector[37] << 3;
assign MEM[301] = input_vector[37] << 2;
assign MEM[302] = input_vector[37] << 1;
assign MEM[303] = input_vector[37] << 0;
assign MEM[304] = -(input_vector[38] << 7);
assign MEM[305] = input_vector[38] << 6;
assign MEM[306] = input_vector[38] << 5;
assign MEM[307] = input_vector[38] << 4;
assign MEM[308] = input_vector[38] << 3;
assign MEM[309] = input_vector[38] << 2;
assign MEM[310] = input_vector[38] << 1;
assign MEM[311] = input_vector[38] << 0;
assign MEM[312] = -(input_vector[39] << 7);
assign MEM[313] = input_vector[39] << 6;
assign MEM[314] = input_vector[39] << 5;
assign MEM[315] = input_vector[39] << 4;
assign MEM[316] = input_vector[39] << 3;
assign MEM[317] = input_vector[39] << 2;
assign MEM[318] = input_vector[39] << 1;
assign MEM[319] = input_vector[39] << 0;
assign MEM[320] = -(input_vector[40] << 7);
assign MEM[321] = input_vector[40] << 6;
assign MEM[322] = input_vector[40] << 5;
assign MEM[323] = input_vector[40] << 4;
assign MEM[324] = input_vector[40] << 3;
assign MEM[325] = input_vector[40] << 2;
assign MEM[326] = input_vector[40] << 1;
assign MEM[327] = input_vector[40] << 0;
assign MEM[328] = -(input_vector[41] << 7);
assign MEM[329] = input_vector[41] << 6;
assign MEM[330] = input_vector[41] << 5;
assign MEM[331] = input_vector[41] << 4;
assign MEM[332] = input_vector[41] << 3;
assign MEM[333] = input_vector[41] << 2;
assign MEM[334] = input_vector[41] << 1;
assign MEM[335] = input_vector[41] << 0;
assign MEM[336] = -(input_vector[42] << 7);
assign MEM[337] = input_vector[42] << 6;
assign MEM[338] = input_vector[42] << 5;
assign MEM[339] = input_vector[42] << 4;
assign MEM[340] = input_vector[42] << 3;
assign MEM[341] = input_vector[42] << 2;
assign MEM[342] = input_vector[42] << 1;
assign MEM[343] = input_vector[42] << 0;
assign MEM[344] = -(input_vector[43] << 7);
assign MEM[345] = input_vector[43] << 6;
assign MEM[346] = input_vector[43] << 5;
assign MEM[347] = input_vector[43] << 4;
assign MEM[348] = input_vector[43] << 3;
assign MEM[349] = input_vector[43] << 2;
assign MEM[350] = input_vector[43] << 1;
assign MEM[351] = input_vector[43] << 0;
assign MEM[352] = -(input_vector[44] << 7);
assign MEM[353] = input_vector[44] << 6;
assign MEM[354] = input_vector[44] << 5;
assign MEM[355] = input_vector[44] << 4;
assign MEM[356] = input_vector[44] << 3;
assign MEM[357] = input_vector[44] << 2;
assign MEM[358] = input_vector[44] << 1;
assign MEM[359] = input_vector[44] << 0;
assign MEM[360] = -(input_vector[45] << 7);
assign MEM[361] = input_vector[45] << 6;
assign MEM[362] = input_vector[45] << 5;
assign MEM[363] = input_vector[45] << 4;
assign MEM[364] = input_vector[45] << 3;
assign MEM[365] = input_vector[45] << 2;
assign MEM[366] = input_vector[45] << 1;
assign MEM[367] = input_vector[45] << 0;
assign MEM[368] = -(input_vector[46] << 7);
assign MEM[369] = input_vector[46] << 6;
assign MEM[370] = input_vector[46] << 5;
assign MEM[371] = input_vector[46] << 4;
assign MEM[372] = input_vector[46] << 3;
assign MEM[373] = input_vector[46] << 2;
assign MEM[374] = input_vector[46] << 1;
assign MEM[375] = input_vector[46] << 0;
assign MEM[376] = -(input_vector[47] << 7);
assign MEM[377] = input_vector[47] << 6;
assign MEM[378] = input_vector[47] << 5;
assign MEM[379] = input_vector[47] << 4;
assign MEM[380] = input_vector[47] << 3;
assign MEM[381] = input_vector[47] << 2;
assign MEM[382] = input_vector[47] << 1;
assign MEM[383] = input_vector[47] << 0;
assign MEM[384] = -(input_vector[48] << 7);
assign MEM[385] = input_vector[48] << 6;
assign MEM[386] = input_vector[48] << 5;
assign MEM[387] = input_vector[48] << 4;
assign MEM[388] = input_vector[48] << 3;
assign MEM[389] = input_vector[48] << 2;
assign MEM[390] = input_vector[48] << 1;
assign MEM[391] = input_vector[48] << 0;
assign MEM[392] = -(input_vector[49] << 7);
assign MEM[393] = input_vector[49] << 6;
assign MEM[394] = input_vector[49] << 5;
assign MEM[395] = input_vector[49] << 4;
assign MEM[396] = input_vector[49] << 3;
assign MEM[397] = input_vector[49] << 2;
assign MEM[398] = input_vector[49] << 1;
assign MEM[399] = input_vector[49] << 0;
assign MEM[400] = -(input_vector[50] << 7);
assign MEM[401] = input_vector[50] << 6;
assign MEM[402] = input_vector[50] << 5;
assign MEM[403] = input_vector[50] << 4;
assign MEM[404] = input_vector[50] << 3;
assign MEM[405] = input_vector[50] << 2;
assign MEM[406] = input_vector[50] << 1;
assign MEM[407] = input_vector[50] << 0;
assign MEM[408] = -(input_vector[51] << 7);
assign MEM[409] = input_vector[51] << 6;
assign MEM[410] = input_vector[51] << 5;
assign MEM[411] = input_vector[51] << 4;
assign MEM[412] = input_vector[51] << 3;
assign MEM[413] = input_vector[51] << 2;
assign MEM[414] = input_vector[51] << 1;
assign MEM[415] = input_vector[51] << 0;
assign MEM[416] = -(input_vector[52] << 7);
assign MEM[417] = input_vector[52] << 6;
assign MEM[418] = input_vector[52] << 5;
assign MEM[419] = input_vector[52] << 4;
assign MEM[420] = input_vector[52] << 3;
assign MEM[421] = input_vector[52] << 2;
assign MEM[422] = input_vector[52] << 1;
assign MEM[423] = input_vector[52] << 0;
assign MEM[424] = -(input_vector[53] << 7);
assign MEM[425] = input_vector[53] << 6;
assign MEM[426] = input_vector[53] << 5;
assign MEM[427] = input_vector[53] << 4;
assign MEM[428] = input_vector[53] << 3;
assign MEM[429] = input_vector[53] << 2;
assign MEM[430] = input_vector[53] << 1;
assign MEM[431] = input_vector[53] << 0;
assign MEM[432] = -(input_vector[54] << 7);
assign MEM[433] = input_vector[54] << 6;
assign MEM[434] = input_vector[54] << 5;
assign MEM[435] = input_vector[54] << 4;
assign MEM[436] = input_vector[54] << 3;
assign MEM[437] = input_vector[54] << 2;
assign MEM[438] = input_vector[54] << 1;
assign MEM[439] = input_vector[54] << 0;
assign MEM[440] = -(input_vector[55] << 7);
assign MEM[441] = input_vector[55] << 6;
assign MEM[442] = input_vector[55] << 5;
assign MEM[443] = input_vector[55] << 4;
assign MEM[444] = input_vector[55] << 3;
assign MEM[445] = input_vector[55] << 2;
assign MEM[446] = input_vector[55] << 1;
assign MEM[447] = input_vector[55] << 0;
assign MEM[448] = -(input_vector[56] << 7);
assign MEM[449] = input_vector[56] << 6;
assign MEM[450] = input_vector[56] << 5;
assign MEM[451] = input_vector[56] << 4;
assign MEM[452] = input_vector[56] << 3;
assign MEM[453] = input_vector[56] << 2;
assign MEM[454] = input_vector[56] << 1;
assign MEM[455] = input_vector[56] << 0;
assign MEM[456] = -(input_vector[57] << 7);
assign MEM[457] = input_vector[57] << 6;
assign MEM[458] = input_vector[57] << 5;
assign MEM[459] = input_vector[57] << 4;
assign MEM[460] = input_vector[57] << 3;
assign MEM[461] = input_vector[57] << 2;
assign MEM[462] = input_vector[57] << 1;
assign MEM[463] = input_vector[57] << 0;
assign MEM[464] = -(input_vector[58] << 7);
assign MEM[465] = input_vector[58] << 6;
assign MEM[466] = input_vector[58] << 5;
assign MEM[467] = input_vector[58] << 4;
assign MEM[468] = input_vector[58] << 3;
assign MEM[469] = input_vector[58] << 2;
assign MEM[470] = input_vector[58] << 1;
assign MEM[471] = input_vector[58] << 0;
assign MEM[472] = -(input_vector[59] << 7);
assign MEM[473] = input_vector[59] << 6;
assign MEM[474] = input_vector[59] << 5;
assign MEM[475] = input_vector[59] << 4;
assign MEM[476] = input_vector[59] << 3;
assign MEM[477] = input_vector[59] << 2;
assign MEM[478] = input_vector[59] << 1;
assign MEM[479] = input_vector[59] << 0;
assign MEM[480] = -(input_vector[60] << 7);
assign MEM[481] = input_vector[60] << 6;
assign MEM[482] = input_vector[60] << 5;
assign MEM[483] = input_vector[60] << 4;
assign MEM[484] = input_vector[60] << 3;
assign MEM[485] = input_vector[60] << 2;
assign MEM[486] = input_vector[60] << 1;
assign MEM[487] = input_vector[60] << 0;
assign MEM[488] = -(input_vector[61] << 7);
assign MEM[489] = input_vector[61] << 6;
assign MEM[490] = input_vector[61] << 5;
assign MEM[491] = input_vector[61] << 4;
assign MEM[492] = input_vector[61] << 3;
assign MEM[493] = input_vector[61] << 2;
assign MEM[494] = input_vector[61] << 1;
assign MEM[495] = input_vector[61] << 0;
assign MEM[496] = -(input_vector[62] << 7);
assign MEM[497] = input_vector[62] << 6;
assign MEM[498] = input_vector[62] << 5;
assign MEM[499] = input_vector[62] << 4;
assign MEM[500] = input_vector[62] << 3;
assign MEM[501] = input_vector[62] << 2;
assign MEM[502] = input_vector[62] << 1;
assign MEM[503] = input_vector[62] << 0;
assign MEM[504] = -(input_vector[63] << 7);
assign MEM[505] = input_vector[63] << 6;
assign MEM[506] = input_vector[63] << 5;
assign MEM[507] = input_vector[63] << 4;
assign MEM[508] = input_vector[63] << 3;
assign MEM[509] = input_vector[63] << 2;
assign MEM[510] = input_vector[63] << 1;
assign MEM[511] = input_vector[63] << 0;
assign MEM[512] = MEM[0] + MEM[488];
assign MEM[513] = MEM[33] + MEM[163];
assign MEM[514] = MEM[171] + MEM[222];
assign MEM[515] = MEM[185] + MEM[357];
assign MEM[516] = MEM[205] + MEM[486];
assign MEM[517] = MEM[216] + MEM[394];
assign MEM[518] = MEM[3] + MEM[48];
assign MEM[519] = MEM[32] + MEM[78];
assign MEM[520] = MEM[162] + MEM[343];
assign MEM[521] = MEM[179] + MEM[513];
assign MEM[522] = MEM[188] + MEM[512];
assign MEM[523] = MEM[217] + MEM[515];
assign MEM[524] = MEM[223] + MEM[277];
assign MEM[525] = MEM[246] + MEM[355];
assign MEM[526] = MEM[287] + MEM[516];
assign MEM[527] = MEM[368] + MEM[524];
assign MEM[528] = MEM[463] + MEM[517];
assign MEM[529] = MEM[514] + MEM[520];
assign MEM[530] = MEM[7] + MEM[269];
assign MEM[531] = MEM[23] + MEM[347];
assign MEM[532] = MEM[34] + MEM[518];
assign MEM[533] = MEM[46] + MEM[264];
assign MEM[534] = MEM[50] + MEM[522];
assign MEM[535] = MEM[54] + MEM[415];
assign MEM[536] = MEM[71] + MEM[184];
assign MEM[537] = MEM[80] + MEM[192];
assign MEM[538] = MEM[112] + MEM[266];
assign MEM[539] = MEM[122] + MEM[442];
assign MEM[540] = MEM[131] + MEM[386];
assign MEM[541] = MEM[139] + MEM[215];
assign MEM[542] = MEM[151] + MEM[160];
assign MEM[543] = MEM[156] + MEM[466];
assign MEM[544] = MEM[172] + MEM[525];
assign MEM[545] = MEM[174] + MEM[284];
assign MEM[546] = MEM[182] + MEM[527];
assign MEM[547] = MEM[193] + MEM[526];
assign MEM[548] = MEM[197] + MEM[296];
assign MEM[549] = MEM[252] + MEM[542];
assign MEM[550] = MEM[262] + MEM[519];
assign MEM[551] = MEM[297] + MEM[523];
assign MEM[552] = MEM[311] + MEM[529];
assign MEM[553] = MEM[324] + MEM[545];
assign MEM[554] = MEM[326] + MEM[521];
assign MEM[555] = MEM[333] + MEM[339];
assign MEM[556] = MEM[358] + MEM[362];
assign MEM[557] = MEM[376] + MEM[377];
assign MEM[558] = MEM[390] + MEM[470];
assign MEM[559] = MEM[502] + MEM[533];
assign MEM[560] = MEM[528] + MEM[532];
assign MEM[561] = MEM[537] + MEM[557];
assign MEM[562] = MEM[538] + MEM[552];
assign MEM[563] = MEM[548] + MEM[551];
assign MEM[564] = MEM[2] + MEM[392];
assign MEM[565] = MEM[15] + MEM[553];
assign MEM[566] = MEM[17] + MEM[265];
assign MEM[567] = MEM[19] + MEM[560];
assign MEM[568] = MEM[28] + MEM[52];
assign MEM[569] = MEM[29] + MEM[484];
assign MEM[570] = MEM[38] + MEM[555];
assign MEM[571] = MEM[39] + MEM[504];
assign MEM[572] = MEM[41] + MEM[541];
assign MEM[573] = MEM[42] + MEM[136];
assign MEM[574] = MEM[47] + MEM[536];
assign MEM[575] = MEM[51] + MEM[340];
assign MEM[576] = MEM[59] + MEM[530];
assign MEM[577] = MEM[67] + MEM[535];
assign MEM[578] = MEM[69] + MEM[198];
assign MEM[579] = MEM[72] + MEM[227];
assign MEM[580] = MEM[75] + MEM[318];
assign MEM[581] = MEM[82] + MEM[261];
assign MEM[582] = MEM[84] + MEM[218];
assign MEM[583] = MEM[85] + MEM[200];
assign MEM[584] = MEM[102] + MEM[366];
assign MEM[585] = MEM[108] + MEM[260];
assign MEM[586] = MEM[109] + MEM[327];
assign MEM[587] = MEM[113] + MEM[491];
assign MEM[588] = MEM[118] + MEM[247];
assign MEM[589] = MEM[130] + MEM[547];
assign MEM[590] = MEM[135] + MEM[539];
assign MEM[591] = MEM[137] + MEM[206];
assign MEM[592] = MEM[146] + MEM[363];
assign MEM[593] = MEM[147] + MEM[173];
assign MEM[594] = MEM[186] + MEM[242];
assign MEM[595] = MEM[203] + MEM[546];
assign MEM[596] = MEM[238] + MEM[534];
assign MEM[597] = MEM[253] + MEM[554];
assign MEM[598] = MEM[274] + MEM[345];
assign MEM[599] = MEM[282] + MEM[370];
assign MEM[600] = MEM[285] + MEM[559];
assign MEM[601] = MEM[291] + MEM[543];
assign MEM[602] = MEM[312] + MEM[313];
assign MEM[603] = MEM[319] + MEM[352];
assign MEM[604] = MEM[328] + MEM[562];
assign MEM[605] = MEM[335] + MEM[544];
assign MEM[606] = MEM[341] + MEM[356];
assign MEM[607] = MEM[342] + MEM[360];
assign MEM[608] = MEM[361] + MEM[540];
assign MEM[609] = MEM[365] + MEM[389];
assign MEM[610] = MEM[378] + MEM[573];
assign MEM[611] = MEM[383] + MEM[578];
assign MEM[612] = MEM[420] + MEM[550];
assign MEM[613] = MEM[439] + MEM[592];
assign MEM[614] = MEM[444] + MEM[531];
assign MEM[615] = MEM[447] + MEM[556];
assign MEM[616] = MEM[453] + MEM[558];
assign MEM[617] = MEM[509] + MEM[569];
assign MEM[618] = MEM[549] + MEM[563];
assign MEM[619] = MEM[580] + MEM[603];
assign MEM[620] = MEM[586] + MEM[616];
assign MEM[621] = MEM[593] + MEM[618];
assign MEM[622] = MEM[598] + MEM[611];
assign MEM[623] = MEM[6] + MEM[49];
assign MEM[624] = MEM[13] + MEM[196];
assign MEM[625] = MEM[16] + MEM[566];
assign MEM[626] = MEM[18] + MEM[571];
assign MEM[627] = MEM[22] + MEM[582];
assign MEM[628] = MEM[24] + MEM[25];
assign MEM[629] = MEM[26] + MEM[37];
assign MEM[630] = MEM[31] + MEM[142];
assign MEM[631] = MEM[40] + MEM[425];
assign MEM[632] = MEM[55] + MEM[338];
assign MEM[633] = MEM[60] + MEM[561];
assign MEM[634] = MEM[62] + MEM[373];
assign MEM[635] = MEM[73] + MEM[306];
assign MEM[636] = MEM[74] + MEM[105];
assign MEM[637] = MEM[77] + MEM[116];
assign MEM[638] = MEM[81] + MEM[201];
assign MEM[639] = MEM[83] + MEM[86];
assign MEM[640] = MEM[87] + MEM[419];
assign MEM[641] = MEM[89] + MEM[350];
assign MEM[642] = MEM[91] + MEM[601];
assign MEM[643] = MEM[92] + MEM[430];
assign MEM[644] = MEM[96] + MEM[612];
assign MEM[645] = MEM[100] + MEM[393];
assign MEM[646] = MEM[101] + MEM[202];
assign MEM[647] = MEM[111] + MEM[213];
assign MEM[648] = MEM[123] + MEM[181];
assign MEM[649] = MEM[127] + MEM[320];
assign MEM[650] = MEM[128] + MEM[290];
assign MEM[651] = MEM[132] + MEM[395];
assign MEM[652] = MEM[141] + MEM[298];
assign MEM[653] = MEM[161] + MEM[602];
assign MEM[654] = MEM[164] + MEM[595];
assign MEM[655] = MEM[166] + MEM[591];
assign MEM[656] = MEM[168] + MEM[396];
assign MEM[657] = MEM[170] + MEM[424];
assign MEM[658] = MEM[176] + MEM[177];
assign MEM[659] = MEM[189] + MEM[388];
assign MEM[660] = MEM[195] + MEM[300];
assign MEM[661] = MEM[204] + MEM[600];
assign MEM[662] = MEM[207] + MEM[594];
assign MEM[663] = MEM[208] + MEM[565];
assign MEM[664] = MEM[210] + MEM[588];
assign MEM[665] = MEM[212] + MEM[351];
assign MEM[666] = MEM[224] + MEM[225];
assign MEM[667] = MEM[226] + MEM[256];
assign MEM[668] = MEM[231] + MEM[332];
assign MEM[669] = MEM[232] + MEM[239];
assign MEM[670] = MEM[237] + MEM[587];
assign MEM[671] = MEM[241] + MEM[570];
assign MEM[672] = MEM[254] + MEM[303];
assign MEM[673] = MEM[257] + MEM[567];
assign MEM[674] = MEM[258] + MEM[613];
assign MEM[675] = MEM[288] + MEM[583];
assign MEM[676] = MEM[292] + MEM[314];
assign MEM[677] = MEM[301] + MEM[622];
assign MEM[678] = MEM[304] + MEM[305];
assign MEM[679] = MEM[307] + MEM[604];
assign MEM[680] = MEM[308] + MEM[346];
assign MEM[681] = MEM[316] + MEM[353];
assign MEM[682] = MEM[321] + MEM[402];
assign MEM[683] = MEM[336] + MEM[391];
assign MEM[684] = MEM[359] + MEM[620];
assign MEM[685] = MEM[369] + MEM[607];
assign MEM[686] = MEM[371] + MEM[596];
assign MEM[687] = MEM[372] + MEM[575];
assign MEM[688] = MEM[375] + MEM[468];
assign MEM[689] = MEM[379] + MEM[615];
assign MEM[690] = MEM[384] + MEM[385];
assign MEM[691] = MEM[401] + MEM[606];
assign MEM[692] = MEM[404] + MEM[508];
assign MEM[693] = MEM[406] + MEM[599];
assign MEM[694] = MEM[408] + MEM[649];
assign MEM[695] = MEM[429] + MEM[585];
assign MEM[696] = MEM[432] + MEM[610];
assign MEM[697] = MEM[433] + MEM[590];
assign MEM[698] = MEM[436] + MEM[660];
assign MEM[699] = MEM[445] + MEM[619];
assign MEM[700] = MEM[450] + MEM[624];
assign MEM[701] = MEM[451] + MEM[576];
assign MEM[702] = MEM[464] + MEM[597];
assign MEM[703] = MEM[472] + MEM[584];
assign MEM[704] = MEM[477] + MEM[617];
assign MEM[705] = MEM[485] + MEM[658];
assign MEM[706] = MEM[494] + MEM[574];
assign MEM[707] = MEM[495] + MEM[577];
assign MEM[708] = MEM[496] + MEM[499];
assign MEM[709] = MEM[498] + MEM[608];
assign MEM[710] = MEM[505] + MEM[506];
assign MEM[711] = MEM[572] + MEM[631];
assign MEM[712] = MEM[579] + MEM[589];
assign MEM[713] = MEM[609] + MEM[621];
assign MEM[714] = MEM[623] + MEM[643];
assign MEM[715] = MEM[628] + MEM[629];
assign MEM[716] = MEM[637] + MEM[650];
assign MEM[717] = MEM[641] + MEM[695];
assign MEM[718] = MEM[647] + MEM[702];
assign MEM[719] = MEM[648] + MEM[677];
assign MEM[720] = MEM[651] + MEM[708];
assign MEM[721] = MEM[665] + MEM[706];
assign MEM[722] = MEM[667] + MEM[673];
assign MEM[723] = MEM[678] + MEM[564];
assign MEM[724] = MEM[680] + MEM[709];
assign MEM[725] = MEM[687] + MEM[581];
assign MEM[726] = MEM[1] + MEM[715];
assign MEM[727] = MEM[14] + MEM[245];
assign MEM[728] = MEM[27] + MEM[614];
assign MEM[729] = MEM[30] + MEM[625];
assign MEM[730] = MEM[36] + MEM[455];
assign MEM[731] = MEM[44] + MEM[657];
assign MEM[732] = MEM[53] + MEM[169];
assign MEM[733] = MEM[56] + MEM[61];
assign MEM[734] = MEM[58] + MEM[299];
assign MEM[735] = MEM[64] + MEM[65];
assign MEM[736] = MEM[66] + MEM[431];
assign MEM[737] = MEM[70] + MEM[692];
assign MEM[738] = MEM[88] + MEM[175];
assign MEM[739] = MEM[93] + MEM[211];
assign MEM[740] = MEM[94] + MEM[190];
assign MEM[741] = MEM[98] + MEM[443];
assign MEM[742] = MEM[99] + MEM[474];
assign MEM[743] = MEM[104] + MEM[302];
assign MEM[744] = MEM[107] + MEM[427];
assign MEM[745] = MEM[110] + MEM[568];
assign MEM[746] = MEM[114] + MEM[120];
assign MEM[747] = MEM[115] + MEM[416];
assign MEM[748] = MEM[121] + MEM[157];
assign MEM[749] = MEM[124] + MEM[150];
assign MEM[750] = MEM[126] + MEM[435];
assign MEM[751] = MEM[129] + MEM[671];
assign MEM[752] = MEM[134] + MEM[138];
assign MEM[753] = MEM[148] + MEM[605];
assign MEM[754] = MEM[153] + MEM[645];
assign MEM[755] = MEM[154] + MEM[315];
assign MEM[756] = MEM[159] + MEM[344];
assign MEM[757] = MEM[187] + MEM[364];
assign MEM[758] = MEM[194] + MEM[639];
assign MEM[759] = MEM[209] + MEM[634];
assign MEM[760] = MEM[220] + MEM[309];
assign MEM[761] = MEM[221] + MEM[418];
assign MEM[762] = MEM[229] + MEM[283];
assign MEM[763] = MEM[233] + MEM[669];
assign MEM[764] = MEM[234] + MEM[635];
assign MEM[765] = MEM[235] + MEM[413];
assign MEM[766] = MEM[236] + MEM[714];
assign MEM[767] = MEM[240] + MEM[662];
assign MEM[768] = MEM[243] + MEM[248];
assign MEM[769] = MEM[249] + MEM[250];
assign MEM[770] = MEM[251] + MEM[686];
assign MEM[771] = MEM[255] + MEM[457];
assign MEM[772] = MEM[263] + MEM[640];
assign MEM[773] = MEM[268] + MEM[638];
assign MEM[774] = MEM[272] + MEM[273];
assign MEM[775] = MEM[278] + MEM[630];
assign MEM[776] = MEM[280] + MEM[654];
assign MEM[777] = MEM[286] + MEM[707];
assign MEM[778] = MEM[294] + MEM[670];
assign MEM[779] = MEM[322] + MEM[428];
assign MEM[780] = MEM[330] + MEM[722];
assign MEM[781] = MEM[337] + MEM[636];
assign MEM[782] = MEM[348] + MEM[467];
assign MEM[783] = MEM[349] + MEM[699];
assign MEM[784] = MEM[367] + MEM[701];
assign MEM[785] = MEM[374] + MEM[652];
assign MEM[786] = MEM[380] + MEM[642];
assign MEM[787] = MEM[381] + MEM[682];
assign MEM[788] = MEM[387] + MEM[476];
assign MEM[789] = MEM[398] + MEM[672];
assign MEM[790] = MEM[400] + MEM[691];
assign MEM[791] = MEM[410] + MEM[492];
assign MEM[792] = MEM[411] + MEM[490];
assign MEM[793] = MEM[414] + MEM[705];
assign MEM[794] = MEM[417] + MEM[685];
assign MEM[795] = MEM[421] + MEM[712];
assign MEM[796] = MEM[434] + MEM[626];
assign MEM[797] = MEM[438] + MEM[710];
assign MEM[798] = MEM[440] + MEM[441];
assign MEM[799] = MEM[452] + MEM[694];
assign MEM[800] = MEM[454] + MEM[655];
assign MEM[801] = MEM[459] + MEM[653];
assign MEM[802] = MEM[473] + MEM[500];
assign MEM[803] = MEM[478] + MEM[679];
assign MEM[804] = MEM[479] + MEM[697];
assign MEM[805] = MEM[480] + MEM[481];
assign MEM[806] = MEM[482] + MEM[761];
assign MEM[807] = MEM[493] + MEM[725];
assign MEM[808] = MEM[497] + MEM[720];
assign MEM[809] = MEM[507] + MEM[719];
assign MEM[810] = MEM[510] + MEM[644];
assign MEM[811] = MEM[511] + MEM[688];
assign MEM[812] = MEM[627] + MEM[656];
assign MEM[813] = MEM[632] + MEM[633];
assign MEM[814] = MEM[646] + MEM[713];
assign MEM[815] = MEM[659] + MEM[675];
assign MEM[816] = MEM[661] + MEM[696];
assign MEM[817] = MEM[663] + MEM[698];
assign MEM[818] = MEM[664] + MEM[668];
assign MEM[819] = MEM[666] + MEM[674];
assign MEM[820] = MEM[676] + MEM[684];
assign MEM[821] = MEM[681] + MEM[700];
assign MEM[822] = MEM[683] + MEM[718];
assign MEM[823] = MEM[689] + MEM[711];
assign MEM[824] = MEM[690] + MEM[721];
assign MEM[825] = MEM[693] + MEM[717];
assign MEM[826] = MEM[703] + MEM[716];
assign MEM[827] = MEM[704] + MEM[745];
assign MEM[828] = MEM[723] + MEM[750];
assign MEM[829] = MEM[732] + MEM[812];
assign MEM[830] = MEM[738] + MEM[825];
assign MEM[831] = MEM[740] + MEM[822];
assign MEM[832] = MEM[743] + MEM[790];
assign MEM[833] = MEM[747] + MEM[794];
assign MEM[834] = MEM[749] + MEM[788];
assign MEM[835] = MEM[756] + MEM[724];
assign MEM[836] = MEM[768] + MEM[769];
assign MEM[837] = MEM[789] + MEM[820];
assign MEM[838] = MEM[805] + MEM[806];
assign MEM[839] = MEM[4] + MEM[437];
assign MEM[840] = MEM[5] + MEM[8];
assign MEM[841] = MEM[9] + MEM[733];
assign MEM[842] = MEM[10] + MEM[731];
assign MEM[843] = MEM[12] + MEM[165];
assign MEM[844] = MEM[20] + MEM[774];
assign MEM[845] = MEM[35] + MEM[178];
assign MEM[846] = MEM[43] + MEM[399];
assign MEM[847] = MEM[57] + MEM[771];
assign MEM[848] = MEM[63] + MEM[751];
assign MEM[849] = MEM[68] + MEM[760];
assign MEM[850] = MEM[90] + MEM[503];
assign MEM[851] = MEM[97] + MEM[469];
assign MEM[852] = MEM[103] + MEM[735];
assign MEM[853] = MEM[106] + MEM[770];
assign MEM[854] = MEM[140] + MEM[730];
assign MEM[855] = MEM[143] + MEM[382];
assign MEM[856] = MEM[149] + MEM[244];
assign MEM[857] = MEM[152] + MEM[471];
assign MEM[858] = MEM[155] + MEM[752];
assign MEM[859] = MEM[167] + MEM[259];
assign MEM[860] = MEM[183] + MEM[739];
assign MEM[861] = MEM[214] + MEM[354];
assign MEM[862] = MEM[228] + MEM[734];
assign MEM[863] = MEM[230] + MEM[736];
assign MEM[864] = MEM[267] + MEM[726];
assign MEM[865] = MEM[271] + MEM[460];
assign MEM[866] = MEM[276] + MEM[289];
assign MEM[867] = MEM[293] + MEM[779];
assign MEM[868] = MEM[295] + MEM[763];
assign MEM[869] = MEM[323] + MEM[334];
assign MEM[870] = MEM[325] + MEM[329];
assign MEM[871] = MEM[331] + MEM[757];
assign MEM[872] = MEM[397] + MEM[817];
assign MEM[873] = MEM[405] + MEM[759];
assign MEM[874] = MEM[407] + MEM[727];
assign MEM[875] = MEM[409] + MEM[799];
assign MEM[876] = MEM[412] + MEM[796];
assign MEM[877] = MEM[426] + MEM[767];
assign MEM[878] = MEM[448] + MEM[449];
assign MEM[879] = MEM[456] + MEM[737];
assign MEM[880] = MEM[458] + MEM[791];
assign MEM[881] = MEM[461] + MEM[729];
assign MEM[882] = MEM[462] + MEM[764];
assign MEM[883] = MEM[465] + MEM[758];
assign MEM[884] = MEM[475] + MEM[787];
assign MEM[885] = MEM[483] + MEM[809];
assign MEM[886] = MEM[489] + MEM[728];
assign MEM[887] = MEM[741] + MEM[793];
assign MEM[888] = MEM[742] + MEM[755];
assign MEM[889] = MEM[744] + MEM[784];
assign MEM[890] = MEM[746] + MEM[748];
assign MEM[891] = MEM[753] + MEM[766];
assign MEM[892] = MEM[754] + MEM[775];
assign MEM[893] = MEM[762] + MEM[776];
assign MEM[894] = MEM[765] + MEM[785];
assign MEM[895] = MEM[772] + MEM[778];
assign MEM[896] = MEM[773] + MEM[781];
assign MEM[897] = MEM[777] + MEM[780];
assign MEM[898] = MEM[782] + MEM[811];
assign MEM[899] = MEM[783] + MEM[792];
assign MEM[900] = MEM[786] + MEM[807];
assign MEM[901] = MEM[797] + MEM[814];
assign MEM[902] = MEM[798] + MEM[802];
assign MEM[903] = MEM[800] + MEM[821];
assign MEM[904] = MEM[801] + MEM[804];
assign MEM[905] = MEM[803] + MEM[826];
assign MEM[906] = MEM[808] + MEM[818];
assign MEM[907] = MEM[810] + MEM[834];
assign MEM[908] = MEM[813] + MEM[830];
assign MEM[909] = MEM[815] + MEM[827];
assign MEM[910] = MEM[816] + MEM[833];
assign MEM[911] = MEM[819] + MEM[845];
assign MEM[912] = MEM[823] + MEM[832];
assign MEM[913] = MEM[828] + MEM[829];
assign MEM[914] = MEM[831] + MEM[836];
assign MEM[915] = MEM[838] + MEM[850];
assign MEM[916] = MEM[841] + MEM[893];
assign MEM[917] = MEM[842] + MEM[903];
assign MEM[918] = MEM[847] + MEM[899];
assign MEM[919] = MEM[852] + MEM[795];
assign MEM[920] = MEM[855] + MEM[906];
assign MEM[921] = MEM[856] + MEM[869];
assign MEM[922] = MEM[857] + MEM[890];
assign MEM[923] = MEM[861] + MEM[886];
assign MEM[924] = MEM[862] + MEM[908];
assign MEM[925] = MEM[865] + MEM[835];
assign MEM[926] = MEM[866] + MEM[877];
assign MEM[927] = MEM[874] + MEM[921];
assign MEM[928] = MEM[878] + MEM[889];
assign MEM[929] = MEM[888] + MEM[911];
assign MEM[930] = MEM[892] + MEM[922];
assign MEM[931] = MEM[897] + MEM[907];
assign MEM[932] = MEM[902] + MEM[905];
assign MEM[933] = MEM[11] + MEM[133];
assign MEM[934] = MEM[21] + MEM[854];
assign MEM[935] = MEM[45] + MEM[849];
assign MEM[936] = MEM[76] + MEM[824];
assign MEM[937] = MEM[79] + MEM[119];
assign MEM[938] = MEM[95] + MEM[423];
assign MEM[939] = MEM[117] + MEM[853];
assign MEM[940] = MEM[125] + MEM[275];
assign MEM[941] = MEM[144] + MEM[145];
assign MEM[942] = MEM[158] + MEM[859];
assign MEM[943] = MEM[180] + MEM[875];
assign MEM[944] = MEM[191] + MEM[270];
assign MEM[945] = MEM[199] + MEM[837];
assign MEM[946] = MEM[219] + MEM[880];
assign MEM[947] = MEM[279] + MEM[840];
assign MEM[948] = MEM[317] + MEM[844];
assign MEM[949] = MEM[403] + MEM[851];
assign MEM[950] = MEM[422] + MEM[879];
assign MEM[951] = MEM[430] + MEM[568];
assign MEM[952] = MEM[446] + MEM[858];
assign MEM[953] = MEM[487] + MEM[860];
assign MEM[954] = MEM[501] + MEM[839];
assign MEM[955] = MEM[561] + MEM[846];
assign MEM[956] = MEM[605] + MEM[872];
assign MEM[957] = MEM[614] + MEM[882];
assign MEM[958] = MEM[824] + MEM[871];
assign MEM[959] = MEM[837] + MEM[873];
assign MEM[960] = MEM[843] + MEM[848];
assign MEM[961] = MEM[863] + MEM[868];
assign MEM[962] = MEM[864] + MEM[867];
assign MEM[963] = MEM[870] + MEM[904];
assign MEM[964] = MEM[876] + MEM[894];
assign MEM[965] = MEM[881] + MEM[891];
assign MEM[966] = MEM[883] + MEM[914];
assign MEM[967] = MEM[884] + MEM[912];
assign MEM[968] = MEM[885] + MEM[887];
assign MEM[969] = MEM[895] + MEM[901];
assign MEM[970] = MEM[896] + MEM[909];
assign MEM[971] = MEM[898] + MEM[931];
assign MEM[972] = MEM[900] + MEM[925];
assign MEM[973] = MEM[910] + MEM[915];
assign MEM[974] = MEM[916] + MEM[918];
assign MEM[975] = MEM[917] + MEM[924];
assign MEM[976] = MEM[919] + MEM[923];
assign MEM[977] = MEM[920] + MEM[932];
assign MEM[978] = MEM[926] + MEM[930];
assign MEM[979] = MEM[927] + MEM[934];
assign MEM[980] = MEM[928] + MEM[936];
assign MEM[981] = MEM[929] + MEM[933];
assign MEM[982] = MEM[935] + MEM[970];
assign MEM[983] = MEM[937] + MEM[951];
assign MEM[984] = MEM[938] + MEM[955];
assign MEM[985] = MEM[942] + MEM[967];
assign MEM[986] = MEM[945] + MEM[960];
assign MEM[987] = MEM[946] + MEM[976];
assign MEM[988] = MEM[948] + MEM[962];
assign MEM[989] = MEM[963] + MEM[978];
assign MEM[990] = MEM[968] + MEM[977];
assign MEM[991] = MEM[969] + MEM[973];
assign MEM[992] = MEM[28] + MEM[49];
assign MEM[993] = MEM[74] + MEM[80];
assign MEM[994] = MEM[82] + MEM[124];
assign MEM[995] = MEM[86] + MEM[226];
assign MEM[996] = MEM[116] + MEM[264];
assign MEM[997] = MEM[120] + MEM[134];
assign MEM[998] = MEM[136] + MEM[202];
assign MEM[999] = MEM[138] + MEM[244];
assign MEM[1000] = MEM[142] + MEM[200];
assign MEM[1001] = MEM[157] + MEM[213];
assign MEM[1002] = MEM[178] + MEM[338];
assign MEM[1003] = MEM[201] + MEM[245];
assign MEM[1004] = MEM[211] + MEM[340];
assign MEM[1005] = MEM[227] + MEM[298];
assign MEM[1006] = MEM[235] + MEM[265];
assign MEM[1007] = MEM[242] + MEM[276];
assign MEM[1008] = MEM[269] + MEM[318];
assign MEM[1009] = MEM[277] + MEM[392];
assign MEM[1010] = MEM[281] + MEM[300];
assign MEM[1011] = MEM[290] + MEM[351];
assign MEM[1012] = MEM[309] + MEM[320];
assign MEM[1013] = MEM[310] + MEM[352];
assign MEM[1014] = MEM[314] + MEM[402];
assign MEM[1015] = MEM[321] + MEM[336];
assign MEM[1016] = MEM[339] + MEM[383];
assign MEM[1017] = MEM[342] + MEM[344];
assign MEM[1018] = MEM[347] + MEM[425];
assign MEM[1019] = MEM[353] + MEM[467];
assign MEM[1020] = MEM[360] + MEM[519];
assign MEM[1021] = MEM[364] + MEM[404];
assign MEM[1022] = MEM[373] + MEM[389];
assign MEM[1023] = MEM[391] + MEM[443];
assign MEM[1024] = MEM[395] + MEM[413];
assign MEM[1025] = MEM[396] + MEM[419];
assign MEM[1026] = MEM[418] + MEM[558];
assign MEM[1027] = MEM[428] + MEM[429];
assign MEM[1028] = MEM[431] + MEM[444];
assign MEM[1029] = MEM[434] + MEM[451];
assign MEM[1030] = MEM[454] + MEM[491];
assign MEM[1031] = MEM[455] + MEM[456];
assign MEM[1032] = MEM[457] + MEM[461];
assign MEM[1033] = MEM[471] + MEM[516];
assign MEM[1034] = MEM[474] + MEM[490];
assign MEM[1035] = MEM[484] + MEM[517];
assign MEM[1036] = MEM[494] + MEM[515];
assign MEM[1037] = MEM[510] + MEM[513];
assign MEM[1038] = MEM[512] + MEM[514];
assign MEM[1039] = MEM[518] + MEM[527];
assign MEM[1040] = MEM[521] + MEM[572];
assign MEM[1041] = MEM[522] + MEM[525];
assign MEM[1042] = MEM[523] + MEM[546];
assign MEM[1043] = MEM[526] + MEM[534];
assign MEM[1044] = MEM[528] + MEM[541];
assign MEM[1045] = MEM[529] + MEM[544];
assign MEM[1046] = MEM[530] + MEM[553];
assign MEM[1047] = MEM[531] + MEM[535];
assign MEM[1048] = MEM[536] + MEM[563];
assign MEM[1049] = MEM[539] + MEM[562];
assign MEM[1050] = MEM[540] + MEM[543];
assign MEM[1051] = MEM[547] + MEM[549];
assign MEM[1052] = MEM[550] + MEM[567];
assign MEM[1053] = MEM[554] + MEM[559];
assign MEM[1054] = MEM[555] + MEM[579];
assign MEM[1055] = MEM[556] + MEM[589];
assign MEM[1056] = MEM[560] + MEM[577];
assign MEM[1057] = MEM[564] + MEM[565];
assign MEM[1058] = MEM[566] + MEM[571];
assign MEM[1059] = MEM[570] + MEM[581];
assign MEM[1060] = MEM[574] + MEM[576];
assign MEM[1061] = MEM[575] + MEM[594];
assign MEM[1062] = MEM[582] + MEM[599];
assign MEM[1063] = MEM[583] + MEM[636];
assign MEM[1064] = MEM[584] + MEM[606];
assign MEM[1065] = MEM[585] + MEM[591];
assign MEM[1066] = MEM[587] + MEM[595];
assign MEM[1067] = MEM[588] + MEM[604];
assign MEM[1068] = MEM[590] + MEM[609];
assign MEM[1069] = MEM[596] + MEM[601];
assign MEM[1070] = MEM[597] + MEM[602];
assign MEM[1071] = MEM[600] + MEM[615];
assign MEM[1072] = MEM[607] + MEM[608];
assign MEM[1073] = MEM[610] + MEM[633];
assign MEM[1074] = MEM[612] + MEM[613];
assign MEM[1075] = MEM[617] + MEM[619];
assign MEM[1076] = MEM[620] + MEM[627];
assign MEM[1077] = MEM[621] + MEM[646];
assign MEM[1078] = MEM[622] + MEM[625];
assign MEM[1079] = MEM[626] + MEM[632];
assign MEM[1080] = MEM[630] + MEM[652];
assign MEM[1081] = MEM[634] + MEM[638];
assign MEM[1082] = MEM[635] + MEM[664];
assign MEM[1083] = MEM[639] + MEM[640];
assign MEM[1084] = MEM[642] + MEM[674];
assign MEM[1085] = MEM[644] + MEM[685];
assign MEM[1086] = MEM[645] + MEM[675];
assign MEM[1087] = MEM[653] + MEM[659];
assign MEM[1088] = MEM[654] + MEM[656];
assign MEM[1089] = MEM[655] + MEM[657];
assign MEM[1090] = MEM[661] + MEM[692];
assign MEM[1091] = MEM[662] + MEM[666];
assign MEM[1092] = MEM[663] + MEM[683];
assign MEM[1093] = MEM[668] + MEM[670];
assign MEM[1094] = MEM[669] + MEM[671];
assign MEM[1095] = MEM[672] + MEM[679];
assign MEM[1096] = MEM[676] + MEM[689];
assign MEM[1097] = MEM[681] + MEM[682];
assign MEM[1098] = MEM[684] + MEM[704];
assign MEM[1099] = MEM[686] + MEM[717];
assign MEM[1100] = MEM[688] + MEM[698];
assign MEM[1101] = MEM[690] + MEM[694];
assign MEM[1102] = MEM[691] + MEM[696];
assign MEM[1103] = MEM[693] + MEM[701];
assign MEM[1104] = MEM[697] + MEM[722];
assign MEM[1105] = MEM[699] + MEM[707];
assign MEM[1106] = MEM[700] + MEM[712];
assign MEM[1107] = MEM[703] + MEM[721];
assign MEM[1108] = MEM[705] + MEM[710];
assign MEM[1109] = MEM[711] + MEM[714];
assign MEM[1110] = MEM[713] + MEM[715];
assign MEM[1111] = MEM[716] + MEM[719];
assign MEM[1112] = MEM[718] + MEM[725];
assign MEM[1113] = MEM[720] + MEM[746];
assign MEM[1114] = MEM[723] + MEM[727];
assign MEM[1115] = MEM[724] + MEM[755];
assign MEM[1116] = MEM[726] + MEM[731];
assign MEM[1117] = MEM[728] + MEM[730];
assign MEM[1118] = MEM[729] + MEM[773];
assign MEM[1119] = MEM[733] + MEM[757];
assign MEM[1120] = MEM[734] + MEM[737];
assign MEM[1121] = MEM[735] + MEM[751];
assign MEM[1122] = MEM[736] + MEM[748];
assign MEM[1123] = MEM[739] + MEM[752];
assign MEM[1124] = MEM[741] + MEM[781];
assign MEM[1125] = MEM[742] + MEM[754];
assign MEM[1126] = MEM[744] + MEM[771];
assign MEM[1127] = MEM[753] + MEM[760];
assign MEM[1128] = MEM[758] + MEM[765];
assign MEM[1129] = MEM[759] + MEM[778];
assign MEM[1130] = MEM[762] + MEM[766];
assign MEM[1131] = MEM[763] + MEM[784];
assign MEM[1132] = MEM[764] + MEM[774];
assign MEM[1133] = MEM[767] + MEM[796];
assign MEM[1134] = MEM[770] + MEM[776];
assign MEM[1135] = MEM[772] + MEM[786];
assign MEM[1136] = MEM[775] + MEM[779];
assign MEM[1137] = MEM[777] + MEM[797];
assign MEM[1138] = MEM[780] + MEM[783];
assign MEM[1139] = MEM[782] + MEM[785];
assign MEM[1140] = MEM[787] + MEM[795];
assign MEM[1141] = MEM[791] + MEM[792];
assign MEM[1142] = MEM[793] + MEM[801];
assign MEM[1143] = MEM[798] + MEM[799];
assign MEM[1144] = MEM[800] + MEM[802];
assign MEM[1145] = MEM[803] + MEM[867];
assign MEM[1146] = MEM[804] + MEM[809];
assign MEM[1147] = MEM[807] + MEM[828];
assign MEM[1148] = MEM[808] + MEM[814];
assign MEM[1149] = MEM[810] + MEM[815];
assign MEM[1150] = MEM[811] + MEM[813];
assign MEM[1151] = MEM[816] + MEM[829];
assign MEM[1152] = MEM[817] + MEM[819];
assign MEM[1153] = MEM[818] + MEM[821];
assign MEM[1154] = MEM[823] + MEM[827];
assign MEM[1155] = MEM[826] + MEM[853];
assign MEM[1156] = MEM[830] + MEM[846];
assign MEM[1157] = MEM[831] + MEM[843];
assign MEM[1158] = MEM[832] + MEM[864];
assign MEM[1159] = MEM[833] + MEM[838];
assign MEM[1160] = MEM[834] + MEM[839];
assign MEM[1161] = MEM[835] + MEM[854];
assign MEM[1162] = MEM[836] + MEM[883];
assign MEM[1163] = MEM[840] + MEM[844];
assign MEM[1164] = MEM[848] + MEM[859];
assign MEM[1165] = MEM[849] + MEM[870];
assign MEM[1166] = MEM[851] + MEM[863];
assign MEM[1167] = MEM[858] + MEM[876];
assign MEM[1168] = MEM[860] + MEM[880];
assign MEM[1169] = MEM[868] + MEM[875];
assign MEM[1170] = MEM[871] + MEM[879];
assign MEM[1171] = MEM[872] + MEM[873];
assign MEM[1172] = MEM[881] + MEM[894];
assign MEM[1173] = MEM[882] + MEM[884];
assign MEM[1174] = MEM[885] + MEM[891];
assign MEM[1175] = MEM[887] + MEM[919];
assign MEM[1176] = MEM[895] + MEM[924];
assign MEM[1177] = MEM[896] + MEM[912];
assign MEM[1178] = MEM[898] + MEM[900];
assign MEM[1179] = MEM[901] + MEM[916];
assign MEM[1180] = MEM[904] + MEM[947];
assign MEM[1181] = MEM[909] + MEM[932];
assign MEM[1182] = MEM[910] + MEM[952];
assign MEM[1183] = MEM[913] + MEM[914];
assign MEM[1184] = MEM[913] + MEM[918];
assign MEM[1185] = MEM[913] + MEM[920];
assign MEM[1186] = MEM[915] + MEM[917];
assign MEM[1187] = MEM[923] + MEM[929];
assign MEM[1188] = MEM[925] + MEM[928];
assign MEM[1189] = MEM[926] + MEM[943];
assign MEM[1190] = MEM[927] + MEM[940];
assign MEM[1191] = MEM[930] + MEM[953];
assign MEM[1192] = MEM[931] + MEM[939];
assign MEM[1193] = MEM[939] + MEM[940];
assign MEM[1194] = MEM[941] + MEM[943];
assign MEM[1195] = MEM[941] + MEM[949];
assign MEM[1196] = MEM[944] + MEM[949];
assign MEM[1197] = MEM[944] + MEM[952];
assign MEM[1198] = MEM[947] + MEM[961];
assign MEM[1199] = MEM[950] + MEM[954];
assign MEM[1200] = MEM[950] + MEM[961];
assign MEM[1201] = MEM[953] + MEM[965];
assign MEM[1202] = MEM[954] + MEM[956];
assign MEM[1203] = MEM[956] + MEM[957];
assign MEM[1204] = MEM[957] + MEM[966];
assign MEM[1205] = MEM[958] + MEM[964];
assign MEM[1206] = MEM[958] + MEM[975];
assign MEM[1207] = MEM[959] + MEM[975];
assign MEM[1208] = MEM[959] + MEM[982];
assign MEM[1209] = MEM[964] + MEM[974];
assign MEM[1210] = MEM[965] + MEM[971];
assign MEM[1211] = MEM[966] + MEM[980];
assign MEM[1212] = MEM[971] + MEM[981];
assign MEM[1213] = MEM[972] + MEM[974];
assign MEM[1214] = MEM[972] + MEM[988];
assign MEM[1215] = MEM[979] + MEM[980];
assign MEM[1216] = MEM[979] + MEM[981];
assign MEM[1217] = MEM[982] + MEM[987];
assign MEM[1218] = MEM[983] + MEM[988];
assign MEM[1219] = MEM[983] + MEM[997];
assign MEM[1220] = MEM[984] + MEM[985];
assign MEM[1221] = MEM[984] + MEM[986];
assign MEM[1222] = MEM[985] + MEM[991];
assign MEM[1223] = MEM[986] + MEM[987];
assign MEM[1224] = MEM[989] + MEM[996];
assign MEM[1225] = MEM[989] + MEM[999];
assign MEM[1226] = MEM[990] + MEM[993];
assign MEM[1227] = MEM[990] + MEM[1005];
assign MEM[1228] = MEM[991] + MEM[1003];
assign MEM[1229] = MEM[992] + MEM[1002];
assign MEM[1230] = MEM[994] + MEM[1006];
assign MEM[1231] = MEM[995] + MEM[1008];
assign MEM[1232] = MEM[998] + MEM[1004];
assign MEM[1233] = MEM[1000] + MEM[1007];
assign MEM[1234] = MEM[1001] + MEM[1014];
assign MEM[1235] = MEM[1009] + MEM[1028];
assign MEM[1236] = MEM[1010] + MEM[1015];
assign MEM[1237] = MEM[1011] + MEM[1025];
assign MEM[1238] = MEM[1012] + MEM[1019];
assign MEM[1239] = MEM[1013] + MEM[1022];
assign MEM[1240] = MEM[1016] + MEM[1024];
assign MEM[1241] = MEM[1017] + MEM[1018];
assign MEM[1242] = MEM[1020] + MEM[1045];
assign MEM[1243] = MEM[1021] + MEM[1026];
assign MEM[1244] = MEM[1023] + MEM[1034];
assign MEM[1245] = MEM[1027] + MEM[1030];
assign MEM[1246] = MEM[1029] + MEM[1031];
assign MEM[1247] = MEM[1032] + MEM[1036];
assign MEM[1248] = MEM[1033] + MEM[1048];
assign MEM[1249] = MEM[1035] + MEM[1041];
assign MEM[1250] = MEM[1037] + MEM[1043];
assign MEM[1251] = MEM[1038] + MEM[1044];
assign MEM[1252] = MEM[1039] + MEM[1058];
assign MEM[1253] = MEM[1040] + MEM[1062];
assign MEM[1254] = MEM[1042] + MEM[1053];
assign MEM[1255] = MEM[1046] + MEM[1055];
assign MEM[1256] = MEM[1047] + MEM[1049];
assign MEM[1257] = MEM[1050] + MEM[1052];
assign MEM[1258] = MEM[1051] + MEM[1054];
assign MEM[1259] = MEM[1056] + MEM[1065];
assign MEM[1260] = MEM[1057] + MEM[1060];
assign MEM[1261] = MEM[1059] + MEM[1068];
assign MEM[1262] = MEM[1061] + MEM[1084];
assign MEM[1263] = MEM[1063] + MEM[1088];
assign MEM[1264] = MEM[1064] + MEM[1082];
assign MEM[1265] = MEM[1066] + MEM[1070];
assign MEM[1266] = MEM[1067] + MEM[1074];
assign MEM[1267] = MEM[1069] + MEM[1073];
assign MEM[1268] = MEM[1071] + MEM[1079];
assign MEM[1269] = MEM[1072] + MEM[1077];
assign MEM[1270] = MEM[1075] + MEM[1078];
assign MEM[1271] = MEM[1076] + MEM[1085];
assign MEM[1272] = MEM[1080] + MEM[1122];
assign MEM[1273] = MEM[1081] + MEM[1098];
assign MEM[1274] = MEM[1083] + MEM[1087];
assign MEM[1275] = MEM[1086] + MEM[1097];
assign MEM[1276] = MEM[1089] + MEM[1093];
assign MEM[1277] = MEM[1090] + MEM[1106];
assign MEM[1278] = MEM[1091] + MEM[1095];
assign MEM[1279] = MEM[1092] + MEM[1099];
assign MEM[1280] = MEM[1094] + MEM[1101];
assign MEM[1281] = MEM[1096] + MEM[1103];
assign MEM[1282] = MEM[1100] + MEM[1105];
assign MEM[1283] = MEM[1102] + MEM[1104];
assign MEM[1284] = MEM[1107] + MEM[1124];
assign MEM[1285] = MEM[1108] + MEM[1109];
assign MEM[1286] = MEM[1110] + MEM[1115];
assign MEM[1287] = MEM[1111] + MEM[1116];
assign MEM[1288] = MEM[1112] + MEM[1118];
assign MEM[1289] = MEM[1113] + MEM[1127];
assign MEM[1290] = MEM[1114] + MEM[1121];
assign MEM[1291] = MEM[1117] + MEM[1126];
assign MEM[1292] = MEM[1119] + MEM[1132];
assign MEM[1293] = MEM[1120] + MEM[1125];
assign MEM[1294] = MEM[1123] + MEM[1130];
assign MEM[1295] = MEM[1128] + MEM[1135];
assign MEM[1296] = MEM[1129] + MEM[1147];
assign MEM[1297] = MEM[1131] + MEM[1146];
assign MEM[1298] = MEM[1133] + MEM[1154];
assign MEM[1299] = MEM[1134] + MEM[1138];
assign MEM[1300] = MEM[1136] + MEM[1139];
assign MEM[1301] = MEM[1137] + MEM[1155];
assign MEM[1302] = MEM[1140] + MEM[1144];
assign MEM[1303] = MEM[1141] + MEM[1143];
assign MEM[1304] = MEM[1142] + MEM[1148];
assign MEM[1305] = MEM[1145] + MEM[1176];
assign MEM[1306] = MEM[1149] + MEM[1157];
assign MEM[1307] = MEM[1150] + MEM[1153];
assign MEM[1308] = MEM[1151] + MEM[1162];
assign MEM[1309] = MEM[1152] + MEM[1158];
assign MEM[1310] = MEM[1156] + MEM[1165];
assign MEM[1311] = MEM[1159] + MEM[1164];
assign MEM[1312] = MEM[1160] + MEM[1163];
assign MEM[1313] = MEM[1161] + MEM[1177];
assign MEM[1314] = MEM[1166] + MEM[1171];
assign MEM[1315] = MEM[1167] + MEM[1174];
assign MEM[1316] = MEM[1168] + MEM[1179];
assign MEM[1317] = MEM[1169] + MEM[1178];
assign MEM[1318] = MEM[1170] + MEM[1172];
assign MEM[1319] = MEM[1173] + MEM[1175];
assign MEM[1320] = MEM[1180] + MEM[1199];
assign MEM[1321] = MEM[1181] + MEM[1195];
assign MEM[1322] = MEM[1182] + MEM[1204];
assign MEM[1323] = MEM[1183] + MEM[1203];
assign MEM[1324] = MEM[1184] + MEM[1189];
assign MEM[1325] = MEM[1185] + MEM[1191];
assign MEM[1326] = MEM[1186] + MEM[1187];
assign MEM[1327] = MEM[1188] + MEM[1198];
assign MEM[1328] = MEM[1190] + MEM[1197];
assign MEM[1329] = MEM[1192] + MEM[1196];
assign MEM[1330] = MEM[1193] + MEM[1194];
assign MEM[1331] = MEM[1200] + MEM[1211];
assign MEM[1332] = MEM[1201] + MEM[1217];
assign MEM[1333] = MEM[1202] + MEM[1214];
assign MEM[1334] = MEM[1205] + MEM[1212];
assign MEM[1335] = MEM[1206] + MEM[1222];
assign MEM[1336] = MEM[1207] + MEM[1215];
assign MEM[1337] = MEM[1208] + MEM[1220];
assign MEM[1338] = MEM[1209] + MEM[1218];
assign MEM[1339] = MEM[1210] + MEM[1226];
assign MEM[1340] = MEM[1213] + MEM[1216];
assign MEM[1341] = MEM[1219] + MEM[1232];
assign MEM[1342] = MEM[1221] + MEM[1225];
assign MEM[1343] = MEM[1223] + MEM[1229];
assign MEM[1344] = MEM[1224] + MEM[1236];
assign MEM[1345] = MEM[1227] + MEM[1239];
assign MEM[1346] = MEM[1228] + MEM[1238];
assign MEM[1347] = MEM[1230] + MEM[1244];
assign MEM[1348] = MEM[1231] + MEM[1240];
assign MEM[1349] = MEM[1233] + MEM[1237];
assign MEM[1350] = MEM[1234] + MEM[1253];
assign MEM[1351] = MEM[1235] + MEM[1255];
assign MEM[1352] = MEM[1241] + MEM[1254];
assign MEM[1353] = MEM[1242] + MEM[1259];
assign MEM[1354] = MEM[1243] + MEM[1260];
assign MEM[1355] = MEM[1245] + MEM[1251];
assign MEM[1356] = MEM[1246] + MEM[1247];
assign MEM[1357] = MEM[1248] + MEM[1265];
assign MEM[1358] = MEM[1249] + MEM[1256];
assign MEM[1359] = MEM[1250] + MEM[1257];
assign MEM[1360] = MEM[1252] + MEM[1266];
assign MEM[1361] = MEM[1258] + MEM[1273];
assign MEM[1362] = MEM[1261] + MEM[1270];
assign MEM[1363] = MEM[1262] + MEM[1281];
assign MEM[1364] = MEM[1263] + MEM[1278];
assign MEM[1365] = MEM[1264] + MEM[1280];
assign MEM[1366] = MEM[1267] + MEM[1275];
assign MEM[1367] = MEM[1268] + MEM[1274];
assign MEM[1368] = MEM[1269] + MEM[1276];
assign MEM[1369] = MEM[1271] + MEM[1283];
assign MEM[1370] = MEM[1272] + MEM[1295];
assign MEM[1371] = MEM[1277] + MEM[1294];
assign MEM[1372] = MEM[1279] + MEM[1293];
assign MEM[1373] = MEM[1282] + MEM[1291];
assign MEM[1374] = MEM[1284] + MEM[1302];
assign MEM[1375] = MEM[1285] + MEM[1288];
assign MEM[1376] = MEM[1286] + MEM[1299];
assign MEM[1377] = MEM[1287] + MEM[1292];
assign MEM[1378] = MEM[1289] + MEM[1297];
assign MEM[1379] = MEM[1290] + MEM[1298];
assign MEM[1380] = MEM[1296] + MEM[1311];
assign MEM[1381] = MEM[1300] + MEM[1304];
assign MEM[1382] = MEM[1301] + MEM[1317];
assign MEM[1383] = MEM[1303] + MEM[1309];
assign MEM[1384] = MEM[1305] + MEM[1328];
assign MEM[1385] = MEM[1306] + MEM[1314];
assign MEM[1386] = MEM[1307] + MEM[1312];
assign MEM[1387] = MEM[1308] + MEM[1321];
assign MEM[1388] = MEM[1310] + MEM[1326];
assign MEM[1389] = MEM[1313] + MEM[1324];
assign MEM[1390] = MEM[1315] + MEM[1320];
assign MEM[1391] = MEM[1316] + MEM[1327];
assign MEM[1392] = MEM[1318] + MEM[1322];
assign MEM[1393] = MEM[1319] + MEM[1329];
assign MEM[1394] = MEM[1323] + MEM[1337];
assign MEM[1395] = MEM[1325] + MEM[1338];
assign MEM[1396] = MEM[1330] + MEM[1333];
assign MEM[1397] = MEM[1331] + MEM[1343];
assign MEM[1398] = MEM[1332] + MEM[1344];
assign MEM[1399] = MEM[1334] + MEM[1342];
assign MEM[1400] = MEM[1335] + MEM[1347];
assign MEM[1401] = MEM[1336] + MEM[1341];
assign MEM[1402] = MEM[1339] + MEM[1350];
assign MEM[1403] = MEM[1340] + MEM[1349];
assign MEM[1404] = MEM[1345] + MEM[1357];
assign MEM[1405] = MEM[1346] + MEM[1358];
assign MEM[1406] = MEM[1348] + MEM[1356];
assign MEM[1407] = MEM[1351] + MEM[1368];
assign MEM[1408] = MEM[1352] + MEM[1362];
assign MEM[1409] = MEM[1353] + MEM[1366];
assign MEM[1410] = MEM[1354] + MEM[1365];
assign MEM[1411] = MEM[1355] + MEM[1361];
assign MEM[1412] = MEM[1359] + MEM[1364];
assign MEM[1413] = MEM[1360] + MEM[1371];
assign MEM[1414] = MEM[1363] + MEM[1374];
assign MEM[1415] = MEM[1367] + MEM[1372];
assign MEM[1416] = MEM[1369] + MEM[1379];
assign MEM[1417] = MEM[1370] + MEM[1383];
assign MEM[1418] = MEM[1373] + MEM[1390];
assign MEM[1419] = MEM[1375] + MEM[1387];
assign MEM[1420] = MEM[1376] + MEM[1384];
assign MEM[1421] = MEM[1377] + MEM[1381];
assign MEM[1422] = MEM[1378] + MEM[1386];
assign MEM[1423] = MEM[1380] + MEM[1391];
assign MEM[1424] = MEM[1382] + MEM[1394];
assign MEM[1425] = MEM[1385] + MEM[1395];
assign MEM[1426] = MEM[1388] + MEM[1396];
assign MEM[1427] = MEM[1389] + MEM[1397];
assign MEM[1428] = MEM[1392] + MEM[1403];
assign MEM[1429] = MEM[1393] + MEM[1401];
assign MEM[1430] = MEM[1398] + MEM[1410];
assign MEM[1431] = MEM[1399] + MEM[1407];
assign MEM[1432] = MEM[1400] + MEM[1412];
assign MEM[1433] = MEM[1402] + MEM[1415];
assign MEM[1434] = MEM[1404] + MEM[1416];
assign MEM[1435] = MEM[1405] + MEM[1414];
assign MEM[1436] = MEM[1406] + MEM[1413];
assign MEM[1437] = MEM[1408] + MEM[1417];
assign MEM[1438] = MEM[1409] + MEM[1421];
assign MEM[1439] = MEM[1411] + MEM[1422];
assign MEM[1440] = MEM[1418] + MEM[1432];
assign MEM[1441] = MEM[1419] + MEM[1431];
assign MEM[1442] = MEM[1420] + MEM[1430];
assign MEM[1443] = MEM[1423] + MEM[1433];
assign MEM[1444] = MEM[1424] + MEM[1436];
assign MEM[1445] = MEM[1425] + MEM[1435];
assign MEM[1446] = MEM[1426] + MEM[1434];
assign MEM[1447] = MEM[1427] + MEM[1438];
assign MEM[1448] = MEM[1428] + MEM[1439];
assign MEM[1449] = MEM[1429] + MEM[1437];
assign output_vector[0] = MEM[1443];
assign output_vector[1] = MEM[1441];
assign output_vector[2] = MEM[1446];
assign output_vector[3] = MEM[1449];
assign output_vector[4] = MEM[1445];
assign output_vector[5] = MEM[1442];
assign output_vector[6] = MEM[1444];
assign output_vector[7] = MEM[1447];
assign output_vector[8] = MEM[1440];
assign output_vector[9] = MEM[1448];

endmodule
