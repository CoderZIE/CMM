// Verilog module
module matrix_mult_optimized_64x64_8_5634#(
    parameter ROWS = 64,
    parameter COLS = 64,
    parameter MEM_SIZE = 5634,
    parameter input_bit_width = 9,
    parameter output_bit_width = 22
)(
    input wire signed [input_bit_width-1:0] input_vector [0: COLS-1],
   output wire signed [output_bit_width-1:0] output_vector [0: ROWS-1]
);

wire signed [output_bit_width-1:0] MEM [0:MEM_SIZE];

assign MEM[0] = -(input_vector[0] << 7);
assign MEM[1] = input_vector[0] << 6;
assign MEM[2] = input_vector[0] << 5;
assign MEM[3] = input_vector[0] << 4;
assign MEM[4] = input_vector[0] << 3;
assign MEM[5] = input_vector[0] << 2;
assign MEM[6] = input_vector[0] << 1;
assign MEM[7] = input_vector[0] << 0;
assign MEM[8] = -(input_vector[1] << 7);
assign MEM[9] = input_vector[1] << 6;
assign MEM[10] = input_vector[1] << 5;
assign MEM[11] = input_vector[1] << 4;
assign MEM[12] = input_vector[1] << 3;
assign MEM[13] = input_vector[1] << 2;
assign MEM[14] = input_vector[1] << 1;
assign MEM[15] = input_vector[1] << 0;
assign MEM[16] = -(input_vector[2] << 7);
assign MEM[17] = input_vector[2] << 6;
assign MEM[18] = input_vector[2] << 5;
assign MEM[19] = input_vector[2] << 4;
assign MEM[20] = input_vector[2] << 3;
assign MEM[21] = input_vector[2] << 2;
assign MEM[22] = input_vector[2] << 1;
assign MEM[23] = input_vector[2] << 0;
assign MEM[24] = -(input_vector[3] << 7);
assign MEM[25] = input_vector[3] << 6;
assign MEM[26] = input_vector[3] << 5;
assign MEM[27] = input_vector[3] << 4;
assign MEM[28] = input_vector[3] << 3;
assign MEM[29] = input_vector[3] << 2;
assign MEM[30] = input_vector[3] << 1;
assign MEM[31] = input_vector[3] << 0;
assign MEM[32] = -(input_vector[4] << 7);
assign MEM[33] = input_vector[4] << 6;
assign MEM[34] = input_vector[4] << 5;
assign MEM[35] = input_vector[4] << 4;
assign MEM[36] = input_vector[4] << 3;
assign MEM[37] = input_vector[4] << 2;
assign MEM[38] = input_vector[4] << 1;
assign MEM[39] = input_vector[4] << 0;
assign MEM[40] = -(input_vector[5] << 7);
assign MEM[41] = input_vector[5] << 6;
assign MEM[42] = input_vector[5] << 5;
assign MEM[43] = input_vector[5] << 4;
assign MEM[44] = input_vector[5] << 3;
assign MEM[45] = input_vector[5] << 2;
assign MEM[46] = input_vector[5] << 1;
assign MEM[47] = input_vector[5] << 0;
assign MEM[48] = -(input_vector[6] << 7);
assign MEM[49] = input_vector[6] << 6;
assign MEM[50] = input_vector[6] << 5;
assign MEM[51] = input_vector[6] << 4;
assign MEM[52] = input_vector[6] << 3;
assign MEM[53] = input_vector[6] << 2;
assign MEM[54] = input_vector[6] << 1;
assign MEM[55] = input_vector[6] << 0;
assign MEM[56] = -(input_vector[7] << 7);
assign MEM[57] = input_vector[7] << 6;
assign MEM[58] = input_vector[7] << 5;
assign MEM[59] = input_vector[7] << 4;
assign MEM[60] = input_vector[7] << 3;
assign MEM[61] = input_vector[7] << 2;
assign MEM[62] = input_vector[7] << 1;
assign MEM[63] = input_vector[7] << 0;
assign MEM[64] = -(input_vector[8] << 7);
assign MEM[65] = input_vector[8] << 6;
assign MEM[66] = input_vector[8] << 5;
assign MEM[67] = input_vector[8] << 4;
assign MEM[68] = input_vector[8] << 3;
assign MEM[69] = input_vector[8] << 2;
assign MEM[70] = input_vector[8] << 1;
assign MEM[71] = input_vector[8] << 0;
assign MEM[72] = -(input_vector[9] << 7);
assign MEM[73] = input_vector[9] << 6;
assign MEM[74] = input_vector[9] << 5;
assign MEM[75] = input_vector[9] << 4;
assign MEM[76] = input_vector[9] << 3;
assign MEM[77] = input_vector[9] << 2;
assign MEM[78] = input_vector[9] << 1;
assign MEM[79] = input_vector[9] << 0;
assign MEM[80] = -(input_vector[10] << 7);
assign MEM[81] = input_vector[10] << 6;
assign MEM[82] = input_vector[10] << 5;
assign MEM[83] = input_vector[10] << 4;
assign MEM[84] = input_vector[10] << 3;
assign MEM[85] = input_vector[10] << 2;
assign MEM[86] = input_vector[10] << 1;
assign MEM[87] = input_vector[10] << 0;
assign MEM[88] = -(input_vector[11] << 7);
assign MEM[89] = input_vector[11] << 6;
assign MEM[90] = input_vector[11] << 5;
assign MEM[91] = input_vector[11] << 4;
assign MEM[92] = input_vector[11] << 3;
assign MEM[93] = input_vector[11] << 2;
assign MEM[94] = input_vector[11] << 1;
assign MEM[95] = input_vector[11] << 0;
assign MEM[96] = -(input_vector[12] << 7);
assign MEM[97] = input_vector[12] << 6;
assign MEM[98] = input_vector[12] << 5;
assign MEM[99] = input_vector[12] << 4;
assign MEM[100] = input_vector[12] << 3;
assign MEM[101] = input_vector[12] << 2;
assign MEM[102] = input_vector[12] << 1;
assign MEM[103] = input_vector[12] << 0;
assign MEM[104] = -(input_vector[13] << 7);
assign MEM[105] = input_vector[13] << 6;
assign MEM[106] = input_vector[13] << 5;
assign MEM[107] = input_vector[13] << 4;
assign MEM[108] = input_vector[13] << 3;
assign MEM[109] = input_vector[13] << 2;
assign MEM[110] = input_vector[13] << 1;
assign MEM[111] = input_vector[13] << 0;
assign MEM[112] = -(input_vector[14] << 7);
assign MEM[113] = input_vector[14] << 6;
assign MEM[114] = input_vector[14] << 5;
assign MEM[115] = input_vector[14] << 4;
assign MEM[116] = input_vector[14] << 3;
assign MEM[117] = input_vector[14] << 2;
assign MEM[118] = input_vector[14] << 1;
assign MEM[119] = input_vector[14] << 0;
assign MEM[120] = -(input_vector[15] << 7);
assign MEM[121] = input_vector[15] << 6;
assign MEM[122] = input_vector[15] << 5;
assign MEM[123] = input_vector[15] << 4;
assign MEM[124] = input_vector[15] << 3;
assign MEM[125] = input_vector[15] << 2;
assign MEM[126] = input_vector[15] << 1;
assign MEM[127] = input_vector[15] << 0;
assign MEM[128] = -(input_vector[16] << 7);
assign MEM[129] = input_vector[16] << 6;
assign MEM[130] = input_vector[16] << 5;
assign MEM[131] = input_vector[16] << 4;
assign MEM[132] = input_vector[16] << 3;
assign MEM[133] = input_vector[16] << 2;
assign MEM[134] = input_vector[16] << 1;
assign MEM[135] = input_vector[16] << 0;
assign MEM[136] = -(input_vector[17] << 7);
assign MEM[137] = input_vector[17] << 6;
assign MEM[138] = input_vector[17] << 5;
assign MEM[139] = input_vector[17] << 4;
assign MEM[140] = input_vector[17] << 3;
assign MEM[141] = input_vector[17] << 2;
assign MEM[142] = input_vector[17] << 1;
assign MEM[143] = input_vector[17] << 0;
assign MEM[144] = -(input_vector[18] << 7);
assign MEM[145] = input_vector[18] << 6;
assign MEM[146] = input_vector[18] << 5;
assign MEM[147] = input_vector[18] << 4;
assign MEM[148] = input_vector[18] << 3;
assign MEM[149] = input_vector[18] << 2;
assign MEM[150] = input_vector[18] << 1;
assign MEM[151] = input_vector[18] << 0;
assign MEM[152] = -(input_vector[19] << 7);
assign MEM[153] = input_vector[19] << 6;
assign MEM[154] = input_vector[19] << 5;
assign MEM[155] = input_vector[19] << 4;
assign MEM[156] = input_vector[19] << 3;
assign MEM[157] = input_vector[19] << 2;
assign MEM[158] = input_vector[19] << 1;
assign MEM[159] = input_vector[19] << 0;
assign MEM[160] = -(input_vector[20] << 7);
assign MEM[161] = input_vector[20] << 6;
assign MEM[162] = input_vector[20] << 5;
assign MEM[163] = input_vector[20] << 4;
assign MEM[164] = input_vector[20] << 3;
assign MEM[165] = input_vector[20] << 2;
assign MEM[166] = input_vector[20] << 1;
assign MEM[167] = input_vector[20] << 0;
assign MEM[168] = -(input_vector[21] << 7);
assign MEM[169] = input_vector[21] << 6;
assign MEM[170] = input_vector[21] << 5;
assign MEM[171] = input_vector[21] << 4;
assign MEM[172] = input_vector[21] << 3;
assign MEM[173] = input_vector[21] << 2;
assign MEM[174] = input_vector[21] << 1;
assign MEM[175] = input_vector[21] << 0;
assign MEM[176] = -(input_vector[22] << 7);
assign MEM[177] = input_vector[22] << 6;
assign MEM[178] = input_vector[22] << 5;
assign MEM[179] = input_vector[22] << 4;
assign MEM[180] = input_vector[22] << 3;
assign MEM[181] = input_vector[22] << 2;
assign MEM[182] = input_vector[22] << 1;
assign MEM[183] = input_vector[22] << 0;
assign MEM[184] = -(input_vector[23] << 7);
assign MEM[185] = input_vector[23] << 6;
assign MEM[186] = input_vector[23] << 5;
assign MEM[187] = input_vector[23] << 4;
assign MEM[188] = input_vector[23] << 3;
assign MEM[189] = input_vector[23] << 2;
assign MEM[190] = input_vector[23] << 1;
assign MEM[191] = input_vector[23] << 0;
assign MEM[192] = -(input_vector[24] << 7);
assign MEM[193] = input_vector[24] << 6;
assign MEM[194] = input_vector[24] << 5;
assign MEM[195] = input_vector[24] << 4;
assign MEM[196] = input_vector[24] << 3;
assign MEM[197] = input_vector[24] << 2;
assign MEM[198] = input_vector[24] << 1;
assign MEM[199] = input_vector[24] << 0;
assign MEM[200] = -(input_vector[25] << 7);
assign MEM[201] = input_vector[25] << 6;
assign MEM[202] = input_vector[25] << 5;
assign MEM[203] = input_vector[25] << 4;
assign MEM[204] = input_vector[25] << 3;
assign MEM[205] = input_vector[25] << 2;
assign MEM[206] = input_vector[25] << 1;
assign MEM[207] = input_vector[25] << 0;
assign MEM[208] = -(input_vector[26] << 7);
assign MEM[209] = input_vector[26] << 6;
assign MEM[210] = input_vector[26] << 5;
assign MEM[211] = input_vector[26] << 4;
assign MEM[212] = input_vector[26] << 3;
assign MEM[213] = input_vector[26] << 2;
assign MEM[214] = input_vector[26] << 1;
assign MEM[215] = input_vector[26] << 0;
assign MEM[216] = -(input_vector[27] << 7);
assign MEM[217] = input_vector[27] << 6;
assign MEM[218] = input_vector[27] << 5;
assign MEM[219] = input_vector[27] << 4;
assign MEM[220] = input_vector[27] << 3;
assign MEM[221] = input_vector[27] << 2;
assign MEM[222] = input_vector[27] << 1;
assign MEM[223] = input_vector[27] << 0;
assign MEM[224] = -(input_vector[28] << 7);
assign MEM[225] = input_vector[28] << 6;
assign MEM[226] = input_vector[28] << 5;
assign MEM[227] = input_vector[28] << 4;
assign MEM[228] = input_vector[28] << 3;
assign MEM[229] = input_vector[28] << 2;
assign MEM[230] = input_vector[28] << 1;
assign MEM[231] = input_vector[28] << 0;
assign MEM[232] = -(input_vector[29] << 7);
assign MEM[233] = input_vector[29] << 6;
assign MEM[234] = input_vector[29] << 5;
assign MEM[235] = input_vector[29] << 4;
assign MEM[236] = input_vector[29] << 3;
assign MEM[237] = input_vector[29] << 2;
assign MEM[238] = input_vector[29] << 1;
assign MEM[239] = input_vector[29] << 0;
assign MEM[240] = -(input_vector[30] << 7);
assign MEM[241] = input_vector[30] << 6;
assign MEM[242] = input_vector[30] << 5;
assign MEM[243] = input_vector[30] << 4;
assign MEM[244] = input_vector[30] << 3;
assign MEM[245] = input_vector[30] << 2;
assign MEM[246] = input_vector[30] << 1;
assign MEM[247] = input_vector[30] << 0;
assign MEM[248] = -(input_vector[31] << 7);
assign MEM[249] = input_vector[31] << 6;
assign MEM[250] = input_vector[31] << 5;
assign MEM[251] = input_vector[31] << 4;
assign MEM[252] = input_vector[31] << 3;
assign MEM[253] = input_vector[31] << 2;
assign MEM[254] = input_vector[31] << 1;
assign MEM[255] = input_vector[31] << 0;
assign MEM[256] = -(input_vector[32] << 7);
assign MEM[257] = input_vector[32] << 6;
assign MEM[258] = input_vector[32] << 5;
assign MEM[259] = input_vector[32] << 4;
assign MEM[260] = input_vector[32] << 3;
assign MEM[261] = input_vector[32] << 2;
assign MEM[262] = input_vector[32] << 1;
assign MEM[263] = input_vector[32] << 0;
assign MEM[264] = -(input_vector[33] << 7);
assign MEM[265] = input_vector[33] << 6;
assign MEM[266] = input_vector[33] << 5;
assign MEM[267] = input_vector[33] << 4;
assign MEM[268] = input_vector[33] << 3;
assign MEM[269] = input_vector[33] << 2;
assign MEM[270] = input_vector[33] << 1;
assign MEM[271] = input_vector[33] << 0;
assign MEM[272] = -(input_vector[34] << 7);
assign MEM[273] = input_vector[34] << 6;
assign MEM[274] = input_vector[34] << 5;
assign MEM[275] = input_vector[34] << 4;
assign MEM[276] = input_vector[34] << 3;
assign MEM[277] = input_vector[34] << 2;
assign MEM[278] = input_vector[34] << 1;
assign MEM[279] = input_vector[34] << 0;
assign MEM[280] = -(input_vector[35] << 7);
assign MEM[281] = input_vector[35] << 6;
assign MEM[282] = input_vector[35] << 5;
assign MEM[283] = input_vector[35] << 4;
assign MEM[284] = input_vector[35] << 3;
assign MEM[285] = input_vector[35] << 2;
assign MEM[286] = input_vector[35] << 1;
assign MEM[287] = input_vector[35] << 0;
assign MEM[288] = -(input_vector[36] << 7);
assign MEM[289] = input_vector[36] << 6;
assign MEM[290] = input_vector[36] << 5;
assign MEM[291] = input_vector[36] << 4;
assign MEM[292] = input_vector[36] << 3;
assign MEM[293] = input_vector[36] << 2;
assign MEM[294] = input_vector[36] << 1;
assign MEM[295] = input_vector[36] << 0;
assign MEM[296] = -(input_vector[37] << 7);
assign MEM[297] = input_vector[37] << 6;
assign MEM[298] = input_vector[37] << 5;
assign MEM[299] = input_vector[37] << 4;
assign MEM[300] = input_vector[37] << 3;
assign MEM[301] = input_vector[37] << 2;
assign MEM[302] = input_vector[37] << 1;
assign MEM[303] = input_vector[37] << 0;
assign MEM[304] = -(input_vector[38] << 7);
assign MEM[305] = input_vector[38] << 6;
assign MEM[306] = input_vector[38] << 5;
assign MEM[307] = input_vector[38] << 4;
assign MEM[308] = input_vector[38] << 3;
assign MEM[309] = input_vector[38] << 2;
assign MEM[310] = input_vector[38] << 1;
assign MEM[311] = input_vector[38] << 0;
assign MEM[312] = -(input_vector[39] << 7);
assign MEM[313] = input_vector[39] << 6;
assign MEM[314] = input_vector[39] << 5;
assign MEM[315] = input_vector[39] << 4;
assign MEM[316] = input_vector[39] << 3;
assign MEM[317] = input_vector[39] << 2;
assign MEM[318] = input_vector[39] << 1;
assign MEM[319] = input_vector[39] << 0;
assign MEM[320] = -(input_vector[40] << 7);
assign MEM[321] = input_vector[40] << 6;
assign MEM[322] = input_vector[40] << 5;
assign MEM[323] = input_vector[40] << 4;
assign MEM[324] = input_vector[40] << 3;
assign MEM[325] = input_vector[40] << 2;
assign MEM[326] = input_vector[40] << 1;
assign MEM[327] = input_vector[40] << 0;
assign MEM[328] = -(input_vector[41] << 7);
assign MEM[329] = input_vector[41] << 6;
assign MEM[330] = input_vector[41] << 5;
assign MEM[331] = input_vector[41] << 4;
assign MEM[332] = input_vector[41] << 3;
assign MEM[333] = input_vector[41] << 2;
assign MEM[334] = input_vector[41] << 1;
assign MEM[335] = input_vector[41] << 0;
assign MEM[336] = -(input_vector[42] << 7);
assign MEM[337] = input_vector[42] << 6;
assign MEM[338] = input_vector[42] << 5;
assign MEM[339] = input_vector[42] << 4;
assign MEM[340] = input_vector[42] << 3;
assign MEM[341] = input_vector[42] << 2;
assign MEM[342] = input_vector[42] << 1;
assign MEM[343] = input_vector[42] << 0;
assign MEM[344] = -(input_vector[43] << 7);
assign MEM[345] = input_vector[43] << 6;
assign MEM[346] = input_vector[43] << 5;
assign MEM[347] = input_vector[43] << 4;
assign MEM[348] = input_vector[43] << 3;
assign MEM[349] = input_vector[43] << 2;
assign MEM[350] = input_vector[43] << 1;
assign MEM[351] = input_vector[43] << 0;
assign MEM[352] = -(input_vector[44] << 7);
assign MEM[353] = input_vector[44] << 6;
assign MEM[354] = input_vector[44] << 5;
assign MEM[355] = input_vector[44] << 4;
assign MEM[356] = input_vector[44] << 3;
assign MEM[357] = input_vector[44] << 2;
assign MEM[358] = input_vector[44] << 1;
assign MEM[359] = input_vector[44] << 0;
assign MEM[360] = -(input_vector[45] << 7);
assign MEM[361] = input_vector[45] << 6;
assign MEM[362] = input_vector[45] << 5;
assign MEM[363] = input_vector[45] << 4;
assign MEM[364] = input_vector[45] << 3;
assign MEM[365] = input_vector[45] << 2;
assign MEM[366] = input_vector[45] << 1;
assign MEM[367] = input_vector[45] << 0;
assign MEM[368] = -(input_vector[46] << 7);
assign MEM[369] = input_vector[46] << 6;
assign MEM[370] = input_vector[46] << 5;
assign MEM[371] = input_vector[46] << 4;
assign MEM[372] = input_vector[46] << 3;
assign MEM[373] = input_vector[46] << 2;
assign MEM[374] = input_vector[46] << 1;
assign MEM[375] = input_vector[46] << 0;
assign MEM[376] = -(input_vector[47] << 7);
assign MEM[377] = input_vector[47] << 6;
assign MEM[378] = input_vector[47] << 5;
assign MEM[379] = input_vector[47] << 4;
assign MEM[380] = input_vector[47] << 3;
assign MEM[381] = input_vector[47] << 2;
assign MEM[382] = input_vector[47] << 1;
assign MEM[383] = input_vector[47] << 0;
assign MEM[384] = -(input_vector[48] << 7);
assign MEM[385] = input_vector[48] << 6;
assign MEM[386] = input_vector[48] << 5;
assign MEM[387] = input_vector[48] << 4;
assign MEM[388] = input_vector[48] << 3;
assign MEM[389] = input_vector[48] << 2;
assign MEM[390] = input_vector[48] << 1;
assign MEM[391] = input_vector[48] << 0;
assign MEM[392] = -(input_vector[49] << 7);
assign MEM[393] = input_vector[49] << 6;
assign MEM[394] = input_vector[49] << 5;
assign MEM[395] = input_vector[49] << 4;
assign MEM[396] = input_vector[49] << 3;
assign MEM[397] = input_vector[49] << 2;
assign MEM[398] = input_vector[49] << 1;
assign MEM[399] = input_vector[49] << 0;
assign MEM[400] = -(input_vector[50] << 7);
assign MEM[401] = input_vector[50] << 6;
assign MEM[402] = input_vector[50] << 5;
assign MEM[403] = input_vector[50] << 4;
assign MEM[404] = input_vector[50] << 3;
assign MEM[405] = input_vector[50] << 2;
assign MEM[406] = input_vector[50] << 1;
assign MEM[407] = input_vector[50] << 0;
assign MEM[408] = -(input_vector[51] << 7);
assign MEM[409] = input_vector[51] << 6;
assign MEM[410] = input_vector[51] << 5;
assign MEM[411] = input_vector[51] << 4;
assign MEM[412] = input_vector[51] << 3;
assign MEM[413] = input_vector[51] << 2;
assign MEM[414] = input_vector[51] << 1;
assign MEM[415] = input_vector[51] << 0;
assign MEM[416] = -(input_vector[52] << 7);
assign MEM[417] = input_vector[52] << 6;
assign MEM[418] = input_vector[52] << 5;
assign MEM[419] = input_vector[52] << 4;
assign MEM[420] = input_vector[52] << 3;
assign MEM[421] = input_vector[52] << 2;
assign MEM[422] = input_vector[52] << 1;
assign MEM[423] = input_vector[52] << 0;
assign MEM[424] = -(input_vector[53] << 7);
assign MEM[425] = input_vector[53] << 6;
assign MEM[426] = input_vector[53] << 5;
assign MEM[427] = input_vector[53] << 4;
assign MEM[428] = input_vector[53] << 3;
assign MEM[429] = input_vector[53] << 2;
assign MEM[430] = input_vector[53] << 1;
assign MEM[431] = input_vector[53] << 0;
assign MEM[432] = -(input_vector[54] << 7);
assign MEM[433] = input_vector[54] << 6;
assign MEM[434] = input_vector[54] << 5;
assign MEM[435] = input_vector[54] << 4;
assign MEM[436] = input_vector[54] << 3;
assign MEM[437] = input_vector[54] << 2;
assign MEM[438] = input_vector[54] << 1;
assign MEM[439] = input_vector[54] << 0;
assign MEM[440] = -(input_vector[55] << 7);
assign MEM[441] = input_vector[55] << 6;
assign MEM[442] = input_vector[55] << 5;
assign MEM[443] = input_vector[55] << 4;
assign MEM[444] = input_vector[55] << 3;
assign MEM[445] = input_vector[55] << 2;
assign MEM[446] = input_vector[55] << 1;
assign MEM[447] = input_vector[55] << 0;
assign MEM[448] = -(input_vector[56] << 7);
assign MEM[449] = input_vector[56] << 6;
assign MEM[450] = input_vector[56] << 5;
assign MEM[451] = input_vector[56] << 4;
assign MEM[452] = input_vector[56] << 3;
assign MEM[453] = input_vector[56] << 2;
assign MEM[454] = input_vector[56] << 1;
assign MEM[455] = input_vector[56] << 0;
assign MEM[456] = -(input_vector[57] << 7);
assign MEM[457] = input_vector[57] << 6;
assign MEM[458] = input_vector[57] << 5;
assign MEM[459] = input_vector[57] << 4;
assign MEM[460] = input_vector[57] << 3;
assign MEM[461] = input_vector[57] << 2;
assign MEM[462] = input_vector[57] << 1;
assign MEM[463] = input_vector[57] << 0;
assign MEM[464] = -(input_vector[58] << 7);
assign MEM[465] = input_vector[58] << 6;
assign MEM[466] = input_vector[58] << 5;
assign MEM[467] = input_vector[58] << 4;
assign MEM[468] = input_vector[58] << 3;
assign MEM[469] = input_vector[58] << 2;
assign MEM[470] = input_vector[58] << 1;
assign MEM[471] = input_vector[58] << 0;
assign MEM[472] = -(input_vector[59] << 7);
assign MEM[473] = input_vector[59] << 6;
assign MEM[474] = input_vector[59] << 5;
assign MEM[475] = input_vector[59] << 4;
assign MEM[476] = input_vector[59] << 3;
assign MEM[477] = input_vector[59] << 2;
assign MEM[478] = input_vector[59] << 1;
assign MEM[479] = input_vector[59] << 0;
assign MEM[480] = -(input_vector[60] << 7);
assign MEM[481] = input_vector[60] << 6;
assign MEM[482] = input_vector[60] << 5;
assign MEM[483] = input_vector[60] << 4;
assign MEM[484] = input_vector[60] << 3;
assign MEM[485] = input_vector[60] << 2;
assign MEM[486] = input_vector[60] << 1;
assign MEM[487] = input_vector[60] << 0;
assign MEM[488] = -(input_vector[61] << 7);
assign MEM[489] = input_vector[61] << 6;
assign MEM[490] = input_vector[61] << 5;
assign MEM[491] = input_vector[61] << 4;
assign MEM[492] = input_vector[61] << 3;
assign MEM[493] = input_vector[61] << 2;
assign MEM[494] = input_vector[61] << 1;
assign MEM[495] = input_vector[61] << 0;
assign MEM[496] = -(input_vector[62] << 7);
assign MEM[497] = input_vector[62] << 6;
assign MEM[498] = input_vector[62] << 5;
assign MEM[499] = input_vector[62] << 4;
assign MEM[500] = input_vector[62] << 3;
assign MEM[501] = input_vector[62] << 2;
assign MEM[502] = input_vector[62] << 1;
assign MEM[503] = input_vector[62] << 0;
assign MEM[504] = -(input_vector[63] << 7);
assign MEM[505] = input_vector[63] << 6;
assign MEM[506] = input_vector[63] << 5;
assign MEM[507] = input_vector[63] << 4;
assign MEM[508] = input_vector[63] << 3;
assign MEM[509] = input_vector[63] << 2;
assign MEM[510] = input_vector[63] << 1;
assign MEM[511] = input_vector[63] << 0;
assign MEM[512] = MEM[280] + MEM[281];
assign MEM[513] = MEM[282] + MEM[512];
assign MEM[514] = MEM[401] + MEM[400];
assign MEM[515] = MEM[224] + MEM[225];
assign MEM[516] = MEM[226] + MEM[515];
assign MEM[517] = MEM[252] + MEM[232];
assign MEM[518] = MEM[488] + MEM[489];
assign MEM[519] = MEM[97] + MEM[96];
assign MEM[520] = MEM[360] + MEM[361];
assign MEM[521] = MEM[120] + MEM[121];
assign MEM[522] = MEM[244] + MEM[75];
assign MEM[523] = MEM[256] + MEM[257];
assign MEM[524] = MEM[298] + MEM[127];
assign MEM[525] = MEM[168] + MEM[169];
assign MEM[526] = MEM[170] + MEM[525];
assign MEM[527] = MEM[337] + MEM[336];
assign MEM[528] = MEM[473] + MEM[472];
assign MEM[529] = MEM[48] + MEM[49];
assign MEM[530] = MEM[193] + MEM[192];
assign MEM[531] = MEM[205] + MEM[37];
assign MEM[532] = MEM[209] + MEM[208];
assign MEM[533] = MEM[236] + MEM[476];
assign MEM[534] = MEM[409] + MEM[408];
assign MEM[535] = MEM[0] + MEM[1];
assign MEM[536] = MEM[24] + MEM[25];
assign MEM[537] = MEM[41] + MEM[40];
assign MEM[538] = MEM[216] + MEM[217];
assign MEM[539] = MEM[233] + MEM[283];
assign MEM[540] = MEM[338] + MEM[61];
assign MEM[541] = MEM[352] + MEM[353];
assign MEM[542] = MEM[372] + MEM[277];
assign MEM[543] = MEM[420] + MEM[188];
assign MEM[544] = MEM[432] + MEM[433];
assign MEM[545] = MEM[9] + MEM[8];
assign MEM[546] = MEM[16] + MEM[17];
assign MEM[547] = MEM[32] + MEM[33];
assign MEM[548] = MEM[50] + MEM[431];
assign MEM[549] = MEM[62] + MEM[331];
assign MEM[550] = MEM[136] + MEM[137];
assign MEM[551] = MEM[234] + MEM[197];
assign MEM[552] = MEM[313] + MEM[312];
assign MEM[553] = MEM[329] + MEM[328];
assign MEM[554] = MEM[513] + MEM[212];
assign MEM[555] = MEM[104] + MEM[105];
assign MEM[556] = MEM[240] + MEM[241];
assign MEM[557] = MEM[248] + MEM[249];
assign MEM[558] = MEM[265] + MEM[264];
assign MEM[559] = MEM[286] + MEM[84];
assign MEM[560] = MEM[303] + MEM[434];
assign MEM[561] = MEM[369] + MEM[368];
assign MEM[562] = MEM[429] + MEM[55];
assign MEM[563] = MEM[450] + MEM[300];
assign MEM[564] = MEM[108] + MEM[7];
assign MEM[565] = MEM[153] + MEM[152];
assign MEM[566] = MEM[187] + MEM[182];
assign MEM[567] = MEM[261] + MEM[46];
assign MEM[568] = MEM[384] + MEM[385];
assign MEM[569] = MEM[423] + MEM[142];
assign MEM[570] = MEM[425] + MEM[424];
assign MEM[571] = MEM[3] + MEM[206];
assign MEM[572] = MEM[23] + MEM[306];
assign MEM[573] = MEM[81] + MEM[80];
assign MEM[574] = MEM[91] + MEM[251];
assign MEM[575] = MEM[94] + MEM[171];
assign MEM[576] = MEM[133] + MEM[98];
assign MEM[577] = MEM[139] + MEM[297];
assign MEM[578] = MEM[147] + MEM[162];
assign MEM[579] = MEM[150] + MEM[214];
assign MEM[580] = MEM[166] + MEM[279];
assign MEM[581] = MEM[167] + MEM[285];
assign MEM[582] = MEM[186] + MEM[254];
assign MEM[583] = MEM[267] + MEM[36];
assign MEM[584] = MEM[296] + MEM[456];
assign MEM[585] = MEM[301] + MEM[27];
assign MEM[586] = MEM[308] + MEM[111];
assign MEM[587] = MEM[310] + MEM[317];
assign MEM[588] = MEM[315] + MEM[148];
assign MEM[589] = MEM[321] + MEM[320];
assign MEM[590] = MEM[323] + MEM[416];
assign MEM[591] = MEM[334] + MEM[191];
assign MEM[592] = MEM[356] + MEM[207];
assign MEM[593] = MEM[393] + MEM[392];
assign MEM[594] = MEM[421] + MEM[441];
assign MEM[595] = MEM[496] + MEM[497];
assign MEM[596] = MEM[29] + MEM[311];
assign MEM[597] = MEM[117] + MEM[278];
assign MEM[598] = MEM[125] + MEM[243];
assign MEM[599] = MEM[129] + MEM[128];
assign MEM[600] = MEM[164] + MEM[179];
assign MEM[601] = MEM[245] + MEM[15];
assign MEM[602] = MEM[276] + MEM[87];
assign MEM[603] = MEM[287] + MEM[382];
assign MEM[604] = MEM[341] + MEM[417];
assign MEM[605] = MEM[366] + MEM[373];
assign MEM[606] = MEM[403] + MEM[146];
assign MEM[607] = MEM[406] + MEM[113];
assign MEM[608] = MEM[410] + MEM[451];
assign MEM[609] = MEM[413] + MEM[457];
assign MEM[610] = MEM[437] + MEM[43];
assign MEM[611] = MEM[462] + MEM[149];
assign MEM[612] = MEM[495] + MEM[260];
assign MEM[613] = MEM[518] + MEM[272];
assign MEM[614] = MEM[12] + MEM[227];
assign MEM[615] = MEM[54] + MEM[343];
assign MEM[616] = MEM[59] + MEM[56];
assign MEM[617] = MEM[72] + MEM[64];
assign MEM[618] = MEM[83] + MEM[238];
assign MEM[619] = MEM[100] + MEM[143];
assign MEM[620] = MEM[103] + MEM[445];
assign MEM[621] = MEM[107] + MEM[381];
assign MEM[622] = MEM[132] + MEM[294];
assign MEM[623] = MEM[134] + MEM[422];
assign MEM[624] = MEM[165] + MEM[430];
assign MEM[625] = MEM[195] + MEM[229];
assign MEM[626] = MEM[215] + MEM[293];
assign MEM[627] = MEM[284] + MEM[349];
assign MEM[628] = MEM[295] + MEM[52];
assign MEM[629] = MEM[326] + MEM[351];
assign MEM[630] = MEM[345] + MEM[344];
assign MEM[631] = MEM[358] + MEM[363];
assign MEM[632] = MEM[376] + MEM[377];
assign MEM[633] = MEM[419] + MEM[258];
assign MEM[634] = MEM[440] + MEM[435];
assign MEM[635] = MEM[482] + MEM[53];
assign MEM[636] = MEM[514] + MEM[39];
assign MEM[637] = MEM[11] + MEM[477];
assign MEM[638] = MEM[18] + MEM[339];
assign MEM[639] = MEM[19] + MEM[402];
assign MEM[640] = MEM[28] + MEM[468];
assign MEM[641] = MEM[31] + MEM[118];
assign MEM[642] = MEM[70] + MEM[516];
assign MEM[643] = MEM[122] + MEM[362];
assign MEM[644] = MEM[126] + MEM[123];
assign MEM[645] = MEM[151] + MEM[469];
assign MEM[646] = MEM[173] + MEM[230];
assign MEM[647] = MEM[178] + MEM[177];
assign MEM[648] = MEM[183] + MEM[228];
assign MEM[649] = MEM[185] + MEM[135];
assign MEM[650] = MEM[200] + MEM[202];
assign MEM[651] = MEM[221] + MEM[268];
assign MEM[652] = MEM[247] + MEM[411];
assign MEM[653] = MEM[253] + MEM[447];
assign MEM[654] = MEM[292] + MEM[379];
assign MEM[655] = MEM[302] + MEM[157];
assign MEM[656] = MEM[389] + MEM[74];
assign MEM[657] = MEM[407] + MEM[428];
assign MEM[658] = MEM[439] + MEM[355];
assign MEM[659] = MEM[448] + MEM[458];
assign MEM[660] = MEM[465] + MEM[395];
assign MEM[661] = MEM[480] + MEM[348];
assign MEM[662] = MEM[483] + MEM[4];
assign MEM[663] = MEM[499] + MEM[180];
assign MEM[664] = MEM[500] + MEM[79];
assign MEM[665] = MEM[510] + MEM[357];
assign MEM[666] = MEM[517] + MEM[269];
assign MEM[667] = MEM[523] + MEM[314];
assign MEM[668] = MEM[647] + MEM[176];
assign MEM[669] = MEM[21] + MEM[342];
assign MEM[670] = MEM[26] + MEM[101];
assign MEM[671] = MEM[44] + MEM[172];
assign MEM[672] = MEM[47] + MEM[262];
assign MEM[673] = MEM[63] + MEM[246];
assign MEM[674] = MEM[65] + MEM[527];
assign MEM[675] = MEM[93] + MEM[196];
assign MEM[676] = MEM[116] + MEM[222];
assign MEM[677] = MEM[141] + MEM[20];
assign MEM[678] = MEM[160] + MEM[340];
assign MEM[679] = MEM[213] + MEM[189];
assign MEM[680] = MEM[218] + MEM[58];
assign MEM[681] = MEM[307] + MEM[82];
assign MEM[682] = MEM[354] + MEM[522];
assign MEM[683] = MEM[370] + MEM[444];
assign MEM[684] = MEM[371] + MEM[492];
assign MEM[685] = MEM[405] + MEM[124];
assign MEM[686] = MEM[470] + MEM[110];
assign MEM[687] = MEM[478] + MEM[42];
assign MEM[688] = MEM[490] + MEM[318];
assign MEM[689] = MEM[504] + MEM[505];
assign MEM[690] = MEM[520] + MEM[521];
assign MEM[691] = MEM[529] + MEM[475];
assign MEM[692] = MEM[38] + MEM[271];
assign MEM[693] = MEM[71] + MEM[275];
assign MEM[694] = MEM[88] + MEM[442];
assign MEM[695] = MEM[112] + MEM[130];
assign MEM[696] = MEM[114] + MEM[364];
assign MEM[697] = MEM[161] + MEM[418];
assign MEM[698] = MEM[184] + MEM[219];
assign MEM[699] = MEM[199] + MEM[386];
assign MEM[700] = MEM[235] + MEM[380];
assign MEM[701] = MEM[291] + MEM[198];
assign MEM[702] = MEM[319] + MEM[95];
assign MEM[703] = MEM[332] + MEM[45];
assign MEM[704] = MEM[335] + MEM[415];
assign MEM[705] = MEM[479] + MEM[305];
assign MEM[706] = MEM[509] + MEM[237];
assign MEM[707] = MEM[511] + MEM[391];
assign MEM[708] = MEM[519] + MEM[5];
assign MEM[709] = MEM[6] + MEM[13];
assign MEM[710] = MEM[35] + MEM[242];
assign MEM[711] = MEM[66] + MEM[76];
assign MEM[712] = MEM[67] + MEM[404];
assign MEM[713] = MEM[68] + MEM[390];
assign MEM[714] = MEM[77] + MEM[346];
assign MEM[715] = MEM[78] + MEM[397];
assign MEM[716] = MEM[86] + MEM[51];
assign MEM[717] = MEM[159] + MEM[73];
assign MEM[718] = MEM[175] + MEM[449];
assign MEM[719] = MEM[201] + MEM[333];
assign MEM[720] = MEM[231] + MEM[464];
assign MEM[721] = MEM[290] + MEM[289];
assign MEM[722] = MEM[322] + MEM[398];
assign MEM[723] = MEM[330] + MEM[115];
assign MEM[724] = MEM[350] + MEM[138];
assign MEM[725] = MEM[367] + MEM[399];
assign MEM[726] = MEM[375] + MEM[526];
assign MEM[727] = MEM[383] + MEM[304];
assign MEM[728] = MEM[394] + MEM[508];
assign MEM[729] = MEM[426] + MEM[436];
assign MEM[730] = MEM[446] + MEM[158];
assign MEM[731] = MEM[481] + MEM[145];
assign MEM[732] = MEM[533] + MEM[466];
assign MEM[733] = MEM[535] + MEM[2];
assign MEM[734] = MEM[538] + MEM[487];
assign MEM[735] = MEM[541] + MEM[544];
assign MEM[736] = MEM[721] + MEM[288];
assign MEM[737] = MEM[724] + MEM[550];
assign MEM[738] = MEM[731] + MEM[144];
assign MEM[739] = MEM[22] + MEM[57];
assign MEM[740] = MEM[69] + MEM[99];
assign MEM[741] = MEM[140] + MEM[388];
assign MEM[742] = MEM[154] + MEM[90];
assign MEM[743] = MEM[155] + MEM[396];
assign MEM[744] = MEM[156] + MEM[455];
assign MEM[745] = MEM[163] + MEM[452];
assign MEM[746] = MEM[210] + MEM[484];
assign MEM[747] = MEM[263] + MEM[553];
assign MEM[748] = MEM[412] + MEM[471];
assign MEM[749] = MEM[414] + MEM[60];
assign MEM[750] = MEM[459] + MEM[498];
assign MEM[751] = MEM[486] + MEM[270];
assign MEM[752] = MEM[494] + MEM[239];
assign MEM[753] = MEM[536] + MEM[325];
assign MEM[754] = MEM[537] + MEM[274];
assign MEM[755] = MEM[539] + MEM[551];
assign MEM[756] = MEM[543] + MEM[443];
assign MEM[757] = MEM[561] + MEM[557];
assign MEM[758] = MEM[89] + MEM[532];
assign MEM[759] = MEM[109] + MEM[531];
assign MEM[760] = MEM[194] + MEM[181];
assign MEM[761] = MEM[204] + MEM[474];
assign MEM[762] = MEM[250] + MEM[131];
assign MEM[763] = MEM[259] + MEM[327];
assign MEM[764] = MEM[299] + MEM[461];
assign MEM[765] = MEM[378] + MEM[540];
assign MEM[766] = MEM[387] + MEM[463];
assign MEM[767] = MEM[485] + MEM[528];
assign MEM[768] = MEM[491] + MEM[534];
assign MEM[769] = MEM[502] + MEM[211];
assign MEM[770] = MEM[524] + MEM[324];
assign MEM[771] = MEM[549] + MEM[562];
assign MEM[772] = MEM[34] + MEM[220];
assign MEM[773] = MEM[92] + MEM[427];
assign MEM[774] = MEM[174] + MEM[546];
assign MEM[775] = MEM[316] + MEM[580];
assign MEM[776] = MEM[347] + MEM[266];
assign MEM[777] = MEM[374] + MEM[14];
assign MEM[778] = MEM[453] + MEM[615];
assign MEM[779] = MEM[501] + MEM[556];
assign MEM[780] = MEM[507] + MEM[506];
assign MEM[781] = MEM[530] + MEM[255];
assign MEM[782] = MEM[542] + MEM[309];
assign MEM[783] = MEM[545] + MEM[555];
assign MEM[784] = MEM[573] + MEM[203];
assign MEM[785] = MEM[10] + MEM[552];
assign MEM[786] = MEM[273] + MEM[547];
assign MEM[787] = MEM[559] + MEM[571];
assign MEM[788] = MEM[563] + MEM[568];
assign MEM[789] = MEM[565] + MEM[570];
assign MEM[790] = MEM[569] + MEM[582];
assign MEM[791] = MEM[589] + MEM[590];
assign MEM[792] = MEM[102] + MEM[566];
assign MEM[793] = MEM[106] + MEM[190];
assign MEM[794] = MEM[119] + MEM[454];
assign MEM[795] = MEM[365] + MEM[503];
assign MEM[796] = MEM[460] + MEM[493];
assign MEM[797] = MEM[548] + MEM[593];
assign MEM[798] = MEM[554] + MEM[558];
assign MEM[799] = MEM[560] + MEM[635];
assign MEM[800] = MEM[564] + MEM[359];
assign MEM[801] = MEM[567] + MEM[85];
assign MEM[802] = MEM[572] + MEM[576];
assign MEM[803] = MEM[581] + MEM[587];
assign MEM[804] = MEM[592] + MEM[591];
assign MEM[805] = MEM[594] + MEM[604];
assign MEM[806] = MEM[599] + MEM[574];
assign MEM[807] = MEM[640] + MEM[613];
assign MEM[808] = MEM[223] + MEM[578];
assign MEM[809] = MEM[438] + MEM[579];
assign MEM[810] = MEM[467] + MEM[597];
assign MEM[811] = MEM[575] + MEM[586];
assign MEM[812] = MEM[577] + MEM[585];
assign MEM[813] = MEM[583] + MEM[675];
assign MEM[814] = MEM[584] + MEM[595];
assign MEM[815] = MEM[596] + MEM[607];
assign MEM[816] = MEM[600] + MEM[625];
assign MEM[817] = MEM[611] + MEM[622];
assign MEM[818] = MEM[617] + MEM[631];
assign MEM[819] = MEM[623] + MEM[643];
assign MEM[820] = MEM[654] + MEM[598];
assign MEM[821] = MEM[659] + MEM[608];
assign MEM[822] = MEM[30] + MEM[605];
assign MEM[823] = MEM[588] + MEM[606];
assign MEM[824] = MEM[601] + MEM[620];
assign MEM[825] = MEM[602] + MEM[651];
assign MEM[826] = MEM[609] + MEM[603];
assign MEM[827] = MEM[610] + MEM[629];
assign MEM[828] = MEM[614] + MEM[633];
assign MEM[829] = MEM[616] + MEM[619];
assign MEM[830] = MEM[618] + MEM[627];
assign MEM[831] = MEM[624] + MEM[672];
assign MEM[832] = MEM[626] + MEM[655];
assign MEM[833] = MEM[632] + MEM[650];
assign MEM[834] = MEM[637] + MEM[661];
assign MEM[835] = MEM[638] + MEM[664];
assign MEM[836] = MEM[648] + MEM[683];
assign MEM[837] = MEM[653] + MEM[684];
assign MEM[838] = MEM[666] + MEM[645];
assign MEM[839] = MEM[688] + MEM[628];
assign MEM[840] = MEM[691] + MEM[649];
assign MEM[841] = MEM[706] + MEM[681];
assign MEM[842] = MEM[727] + MEM[644];
assign MEM[843] = MEM[612] + MEM[621];
assign MEM[844] = MEM[630] + MEM[347];
assign MEM[845] = MEM[636] + MEM[639];
assign MEM[846] = MEM[641] + MEM[317];
assign MEM[847] = MEM[642] + MEM[656];
assign MEM[848] = MEM[646] + MEM[668];
assign MEM[849] = MEM[652] + MEM[658];
assign MEM[850] = MEM[660] + MEM[663];
assign MEM[851] = MEM[662] + MEM[685];
assign MEM[852] = MEM[679] + MEM[680];
assign MEM[853] = MEM[689] + MEM[701];
assign MEM[854] = MEM[702] + MEM[634];
assign MEM[855] = MEM[735] + MEM[677];
assign MEM[856] = MEM[657] + MEM[491];
assign MEM[857] = MEM[665] + MEM[447];
assign MEM[858] = MEM[667] + MEM[534];
assign MEM[859] = MEM[669] + MEM[417];
assign MEM[860] = MEM[670] + MEM[690];
assign MEM[861] = MEM[673] + MEM[687];
assign MEM[862] = MEM[674] + MEM[273];
assign MEM[863] = MEM[676] + MEM[711];
assign MEM[864] = MEM[678] + MEM[276];
assign MEM[865] = MEM[682] + MEM[194];
assign MEM[866] = MEM[686] + MEM[507];
assign MEM[867] = MEM[693] + MEM[694];
assign MEM[868] = MEM[695] + MEM[696];
assign MEM[869] = MEM[698] + MEM[738];
assign MEM[870] = MEM[703] + MEM[699];
assign MEM[871] = MEM[704] + MEM[720];
assign MEM[872] = MEM[707] + MEM[730];
assign MEM[873] = MEM[708] + MEM[722];
assign MEM[874] = MEM[712] + MEM[743];
assign MEM[875] = MEM[723] + MEM[725];
assign MEM[876] = MEM[744] + MEM[728];
assign MEM[877] = MEM[757] + MEM[751];
assign MEM[878] = MEM[205] + MEM[315];
assign MEM[879] = MEM[547] + MEM[710];
assign MEM[880] = MEM[671] + MEM[524];
assign MEM[881] = MEM[692] + MEM[513];
assign MEM[882] = MEM[697] + MEM[419];
assign MEM[883] = MEM[700] + MEM[714];
assign MEM[884] = MEM[705] + MEM[254];
assign MEM[885] = MEM[713] + MEM[746];
assign MEM[886] = MEM[715] + MEM[745];
assign MEM[887] = MEM[716] + MEM[179];
assign MEM[888] = MEM[719] + MEM[750];
assign MEM[889] = MEM[726] + MEM[438];
assign MEM[890] = MEM[733] + MEM[761];
assign MEM[891] = MEM[734] + MEM[77];
assign MEM[892] = MEM[736] + MEM[764];
assign MEM[893] = MEM[737] + MEM[509];
assign MEM[894] = MEM[742] + MEM[71];
assign MEM[895] = MEM[754] + MEM[717];
assign MEM[896] = MEM[778] + MEM[383];
assign MEM[897] = MEM[13] + MEM[233];
assign MEM[898] = MEM[26] + MEM[560];
assign MEM[899] = MEM[68] + MEM[598];
assign MEM[900] = MEM[92] + MEM[681];
assign MEM[901] = MEM[98] + MEM[739];
assign MEM[902] = MEM[111] + MEM[493];
assign MEM[903] = MEM[119] + MEM[709];
assign MEM[904] = MEM[131] + MEM[729];
assign MEM[905] = MEM[139] + MEM[774];
assign MEM[906] = MEM[183] + MEM[108];
assign MEM[907] = MEM[187] + MEM[150];
assign MEM[908] = MEM[196] + MEM[309];
assign MEM[909] = MEM[201] + MEM[310];
assign MEM[910] = MEM[239] + MEM[478];
assign MEM[911] = MEM[245] + MEM[766];
assign MEM[912] = MEM[266] + MEM[756];
assign MEM[913] = MEM[279] + MEM[140];
assign MEM[914] = MEM[295] + MEM[718];
assign MEM[915] = MEM[316] + MEM[596];
assign MEM[916] = MEM[404] + MEM[753];
assign MEM[917] = MEM[420] + MEM[678];
assign MEM[918] = MEM[422] + MEM[100];
assign MEM[919] = MEM[427] + MEM[439];
assign MEM[920] = MEM[431] + MEM[195];
assign MEM[921] = MEM[450] + MEM[151];
assign MEM[922] = MEM[456] + MEM[784];
assign MEM[923] = MEM[461] + MEM[161];
assign MEM[924] = MEM[467] + MEM[519];
assign MEM[925] = MEM[482] + MEM[541];
assign MEM[926] = MEM[502] + MEM[740];
assign MEM[927] = MEM[508] + MEM[284];
assign MEM[928] = MEM[520] + MEM[362];
assign MEM[929] = MEM[528] + MEM[59];
assign MEM[930] = MEM[530] + MEM[142];
assign MEM[931] = MEM[546] + MEM[759];
assign MEM[932] = MEM[554] + MEM[749];
assign MEM[933] = MEM[632] + MEM[603];
assign MEM[934] = MEM[652] + MEM[28];
assign MEM[935] = MEM[732] + MEM[671];
assign MEM[936] = MEM[741] + MEM[178];
assign MEM[937] = MEM[747] + MEM[406];
assign MEM[938] = MEM[748] + MEM[69];
assign MEM[939] = MEM[752] + MEM[62];
assign MEM[940] = MEM[755] + MEM[38];
assign MEM[941] = MEM[758] + MEM[210];
assign MEM[942] = MEM[760] + MEM[578];
assign MEM[943] = MEM[763] + MEM[783];
assign MEM[944] = MEM[765] + MEM[434];
assign MEM[945] = MEM[769] + MEM[396];
assign MEM[946] = MEM[770] + MEM[767];
assign MEM[947] = MEM[771] + MEM[190];
assign MEM[948] = MEM[772] + MEM[126];
assign MEM[949] = MEM[776] + MEM[540];
assign MEM[950] = MEM[777] + MEM[213];
assign MEM[951] = MEM[780] + MEM[389];
assign MEM[952] = MEM[781] + MEM[10];
assign MEM[953] = MEM[785] + MEM[12];
assign MEM[954] = MEM[789] + MEM[99];
assign MEM[955] = MEM[791] + MEM[20];
assign MEM[956] = MEM[5] + MEM[296];
assign MEM[957] = MEM[6] + MEM[102];
assign MEM[958] = MEM[7] + MEM[620];
assign MEM[959] = MEM[15] + MEM[570];
assign MEM[960] = MEM[19] + MEM[22];
assign MEM[961] = MEM[21] + MEM[382];
assign MEM[962] = MEM[29] + MEM[798];
assign MEM[963] = MEM[35] + MEM[371];
assign MEM[964] = MEM[42] + MEM[148];
assign MEM[965] = MEM[43] + MEM[116];
assign MEM[966] = MEM[51] + MEM[314];
assign MEM[967] = MEM[54] + MEM[143];
assign MEM[968] = MEM[57] + MEM[602];
assign MEM[969] = MEM[67] + MEM[236];
assign MEM[970] = MEM[74] + MEM[510];
assign MEM[971] = MEM[78] + MEM[607];
assign MEM[972] = MEM[83] + MEM[773];
assign MEM[973] = MEM[86] + MEM[94];
assign MEM[974] = MEM[101] + MEM[548];
assign MEM[975] = MEM[103] + MEM[327];
assign MEM[976] = MEM[107] + MEM[356];
assign MEM[977] = MEM[122] + MEM[386];
assign MEM[978] = MEM[124] + MEM[159];
assign MEM[979] = MEM[127] + MEM[481];
assign MEM[980] = MEM[132] + MEM[782];
assign MEM[981] = MEM[133] + MEM[167];
assign MEM[982] = MEM[156] + MEM[470];
assign MEM[983] = MEM[162] + MEM[301];
assign MEM[984] = MEM[163] + MEM[275];
assign MEM[985] = MEM[164] + MEM[218];
assign MEM[986] = MEM[165] + MEM[333];
assign MEM[987] = MEM[166] + MEM[14];
assign MEM[988] = MEM[173] + MEM[372];
assign MEM[989] = MEM[177] + MEM[244];
assign MEM[990] = MEM[184] + MEM[185];
assign MEM[991] = MEM[184] + MEM[792];
assign MEM[992] = MEM[189] + MEM[308];
assign MEM[993] = MEM[197] + MEM[3];
assign MEM[994] = MEM[199] + MEM[106];
assign MEM[995] = MEM[211] + MEM[402];
assign MEM[996] = MEM[212] + MEM[517];
assign MEM[997] = MEM[214] + MEM[413];
assign MEM[998] = MEM[221] + MEM[39];
assign MEM[999] = MEM[231] + MEM[436];
assign MEM[1000] = MEM[234] + MEM[593];
assign MEM[1001] = MEM[235] + MEM[452];
assign MEM[1002] = MEM[237] + MEM[805];
assign MEM[1003] = MEM[242] + MEM[516];
assign MEM[1004] = MEM[243] + MEM[503];
assign MEM[1005] = MEM[253] + MEM[160];
assign MEM[1006] = MEM[255] + MEM[198];
assign MEM[1007] = MEM[259] + MEM[480];
assign MEM[1008] = MEM[261] + MEM[796];
assign MEM[1009] = MEM[267] + MEM[468];
assign MEM[1010] = MEM[268] + MEM[412];
assign MEM[1011] = MEM[294] + MEM[559];
assign MEM[1012] = MEM[298] + MEM[307];
assign MEM[1013] = MEM[304] + MEM[572];
assign MEM[1014] = MEM[318] + MEM[500];
assign MEM[1015] = MEM[319] + MEM[762];
assign MEM[1016] = MEM[322] + MEM[445];
assign MEM[1017] = MEM[323] + MEM[341];
assign MEM[1018] = MEM[325] + MEM[394];
assign MEM[1019] = MEM[334] + MEM[600];
assign MEM[1020] = MEM[339] + MEM[552];
assign MEM[1021] = MEM[343] + MEM[381];
assign MEM[1022] = MEM[346] + MEM[611];
assign MEM[1023] = MEM[354] + MEM[365];
assign MEM[1024] = MEM[375] + MEM[418];
assign MEM[1025] = MEM[378] + MEM[484];
assign MEM[1026] = MEM[379] + MEM[459];
assign MEM[1027] = MEM[391] + MEM[466];
assign MEM[1028] = MEM[398] + MEM[775];
assign MEM[1029] = MEM[415] + MEM[588];
assign MEM[1030] = MEM[423] + MEM[297];
assign MEM[1031] = MEM[446] + MEM[621];
assign MEM[1032] = MEM[449] + MEM[172];
assign MEM[1033] = MEM[453] + MEM[395];
assign MEM[1034] = MEM[454] + MEM[665];
assign MEM[1035] = MEM[458] + MEM[410];
assign MEM[1036] = MEM[460] + MEM[538];
assign MEM[1037] = MEM[462] + MEM[387];
assign MEM[1038] = MEM[463] + MEM[324];
assign MEM[1039] = MEM[474] + MEM[630];
assign MEM[1040] = MEM[479] + MEM[657];
assign MEM[1041] = MEM[483] + MEM[511];
assign MEM[1042] = MEM[487] + MEM[428];
assign MEM[1043] = MEM[499] + MEM[601];
assign MEM[1044] = MEM[531] + MEM[605];
assign MEM[1045] = MEM[532] + MEM[690];
assign MEM[1046] = MEM[558] + MEM[631];
assign MEM[1047] = MEM[562] + MEM[348];
assign MEM[1048] = MEM[577] + MEM[706];
assign MEM[1049] = MEM[583] + MEM[358];
assign MEM[1050] = MEM[584] + MEM[171];
assign MEM[1051] = MEM[626] + MEM[46];
assign MEM[1052] = MEM[636] + MEM[779];
assign MEM[1053] = MEM[639] + MEM[287];
assign MEM[1054] = MEM[656] + MEM[725];
assign MEM[1055] = MEM[693] + MEM[713];
assign MEM[1056] = MEM[756] + MEM[291];
assign MEM[1057] = MEM[768] + MEM[223];
assign MEM[1058] = MEM[787] + MEM[569];
assign MEM[1059] = MEM[788] + MEM[421];
assign MEM[1060] = MEM[790] + MEM[263];
assign MEM[1061] = MEM[795] + MEM[634];
assign MEM[1062] = MEM[797] + MEM[627];
assign MEM[1063] = MEM[802] + MEM[262];
assign MEM[1064] = MEM[807] + MEM[663];
assign MEM[1065] = MEM[809] + MEM[335];
assign MEM[1066] = MEM[811] + MEM[93];
assign MEM[1067] = MEM[813] + MEM[542];
assign MEM[1068] = MEM[828] + MEM[357];
assign MEM[1069] = MEM[830] + MEM[31];
assign MEM[1070] = MEM[11] + MEM[18];
assign MEM[1071] = MEM[23] + MEM[182];
assign MEM[1072] = MEM[27] + MEM[407];
assign MEM[1073] = MEM[30] + MEM[61];
assign MEM[1074] = MEM[34] + MEM[574];
assign MEM[1075] = MEM[44] + MEM[110];
assign MEM[1076] = MEM[45] + MEM[70];
assign MEM[1077] = MEM[47] + MEM[543];
assign MEM[1078] = MEM[50] + MEM[390];
assign MEM[1079] = MEM[52] + MEM[130];
assign MEM[1080] = MEM[55] + MEM[277];
assign MEM[1081] = MEM[58] + MEM[283];
assign MEM[1082] = MEM[60] + MEM[330];
assign MEM[1083] = MEM[63] + MEM[556];
assign MEM[1084] = MEM[65] + MEM[403];
assign MEM[1085] = MEM[66] + MEM[149];
assign MEM[1086] = MEM[73] + MEM[522];
assign MEM[1087] = MEM[75] + MEM[230];
assign MEM[1088] = MEM[76] + MEM[141];
assign MEM[1089] = MEM[79] + MEM[364];
assign MEM[1090] = MEM[84] + MEM[200];
assign MEM[1091] = MEM[85] + MEM[568];
assign MEM[1092] = MEM[87] + MEM[688];
assign MEM[1093] = MEM[88] + MEM[521];
assign MEM[1094] = MEM[91] + MEM[526];
assign MEM[1095] = MEM[95] + MEM[270];
assign MEM[1096] = MEM[109] + MEM[485];
assign MEM[1097] = MEM[112] + MEM[388];
assign MEM[1098] = MEM[114] + MEM[645];
assign MEM[1099] = MEM[117] + MEM[191];
assign MEM[1100] = MEM[118] + MEM[292];
assign MEM[1101] = MEM[123] + MEM[299];
assign MEM[1102] = MEM[125] + MEM[286];
assign MEM[1103] = MEM[135] + MEM[158];
assign MEM[1104] = MEM[139] + MEM[529];
assign MEM[1105] = MEM[147] + MEM[545];
assign MEM[1106] = MEM[155] + MEM[146];
assign MEM[1107] = MEM[159] + MEM[247];
assign MEM[1108] = MEM[164] + MEM[820];
assign MEM[1109] = MEM[174] + MEM[250];
assign MEM[1110] = MEM[175] + MEM[614];
assign MEM[1111] = MEM[180] + MEM[238];
assign MEM[1112] = MEM[186] + MEM[719];
assign MEM[1113] = MEM[202] + MEM[205];
assign MEM[1114] = MEM[203] + MEM[707];
assign MEM[1115] = MEM[206] + MEM[477];
assign MEM[1116] = MEM[220] + MEM[405];
assign MEM[1117] = MEM[227] + MEM[303];
assign MEM[1118] = MEM[228] + MEM[687];
assign MEM[1119] = MEM[240] + MEM[134];
assign MEM[1120] = MEM[246] + MEM[498];
assign MEM[1121] = MEM[252] + MEM[293];
assign MEM[1122] = MEM[258] + MEM[533];
assign MEM[1123] = MEM[260] + MEM[102];
assign MEM[1124] = MEM[269] + MEM[815];
assign MEM[1125] = MEM[271] + MEM[698];
assign MEM[1126] = MEM[278] + MEM[490];
assign MEM[1127] = MEM[285] + MEM[443];
assign MEM[1128] = MEM[290] + MEM[827];
assign MEM[1129] = MEM[305] + MEM[338];
assign MEM[1130] = MEM[311] + MEM[332];
assign MEM[1131] = MEM[326] + MEM[549];
assign MEM[1132] = MEM[349] + MEM[604];
assign MEM[1133] = MEM[351] + MEM[591];
assign MEM[1134] = MEM[366] + MEM[705];
assign MEM[1135] = MEM[374] + MEM[440];
assign MEM[1136] = MEM[380] + MEM[426];
assign MEM[1137] = MEM[397] + MEM[595];
assign MEM[1138] = MEM[399] + MEM[544];
assign MEM[1139] = MEM[405] + MEM[435];
assign MEM[1140] = MEM[411] + MEM[299];
assign MEM[1141] = MEM[414] + MEM[430];
assign MEM[1142] = MEM[416] + MEM[799];
assign MEM[1143] = MEM[429] + MEM[448];
assign MEM[1144] = MEM[437] + MEM[486];
assign MEM[1145] = MEM[441] + MEM[609];
assign MEM[1146] = MEM[442] + MEM[539];
assign MEM[1147] = MEM[444] + MEM[668];
assign MEM[1148] = MEM[455] + MEM[571];
assign MEM[1149] = MEM[457] + MEM[469];
assign MEM[1150] = MEM[462] + MEM[567];
assign MEM[1151] = MEM[471] + MEM[674];
assign MEM[1152] = MEM[471] + MEM[722];
assign MEM[1153] = MEM[475] + MEM[649];
assign MEM[1154] = MEM[476] + MEM[612];
assign MEM[1155] = MEM[492] + MEM[610];
assign MEM[1156] = MEM[494] + MEM[518];
assign MEM[1157] = MEM[501] + MEM[566];
assign MEM[1158] = MEM[510] + MEM[643];
assign MEM[1159] = MEM[514] + MEM[54];
assign MEM[1160] = MEM[536] + MEM[606];
assign MEM[1161] = MEM[537] + MEM[786];
assign MEM[1162] = MEM[553] + MEM[215];
assign MEM[1163] = MEM[555] + MEM[552];
assign MEM[1164] = MEM[563] + MEM[629];
assign MEM[1165] = MEM[564] + MEM[422];
assign MEM[1166] = MEM[575] + MEM[658];
assign MEM[1167] = MEM[576] + MEM[793];
assign MEM[1168] = MEM[579] + MEM[646];
assign MEM[1169] = MEM[580] + MEM[670];
assign MEM[1170] = MEM[581] + MEM[740];
assign MEM[1171] = MEM[585] + MEM[565];
assign MEM[1172] = MEM[586] + MEM[729];
assign MEM[1173] = MEM[587] + MEM[669];
assign MEM[1174] = MEM[590] + MEM[865];
assign MEM[1175] = MEM[592] + MEM[825];
assign MEM[1176] = MEM[594] + MEM[728];
assign MEM[1177] = MEM[597] + MEM[801];
assign MEM[1178] = MEM[608] + MEM[637];
assign MEM[1179] = MEM[613] + MEM[619];
assign MEM[1180] = MEM[616] + MEM[680];
assign MEM[1181] = MEM[617] + MEM[804];
assign MEM[1182] = MEM[618] + MEM[502];
assign MEM[1183] = MEM[624] + MEM[82];
assign MEM[1184] = MEM[628] + MEM[697];
assign MEM[1185] = MEM[633] + MEM[499];
assign MEM[1186] = MEM[638] + MEM[524];
assign MEM[1187] = MEM[642] + MEM[676];
assign MEM[1188] = MEM[648] + MEM[835];
assign MEM[1189] = MEM[651] + MEM[300];
assign MEM[1190] = MEM[661] + MEM[686];
assign MEM[1191] = MEM[666] + MEM[768];
assign MEM[1192] = MEM[682] + MEM[232];
assign MEM[1193] = MEM[685] + MEM[561];
assign MEM[1194] = MEM[692] + MEM[747];
assign MEM[1195] = MEM[694] + MEM[736];
assign MEM[1196] = MEM[700] + MEM[285];
assign MEM[1197] = MEM[701] + MEM[662];
assign MEM[1198] = MEM[704] + MEM[609];
assign MEM[1199] = MEM[709] + MEM[495];
assign MEM[1200] = MEM[714] + MEM[500];
assign MEM[1201] = MEM[735] + MEM[691];
assign MEM[1202] = MEM[737] + MEM[573];
assign MEM[1203] = MEM[739] + MEM[166];
assign MEM[1204] = MEM[752] + MEM[803];
assign MEM[1205] = MEM[767] + MEM[708];
assign MEM[1206] = MEM[784] + MEM[644];
assign MEM[1207] = MEM[794] + MEM[23];
assign MEM[1208] = MEM[800] + MEM[817];
assign MEM[1209] = MEM[806] + MEM[89];
assign MEM[1210] = MEM[812] + MEM[846];
assign MEM[1211] = MEM[814] + MEM[536];
assign MEM[1212] = MEM[816] + MEM[207];
assign MEM[1213] = MEM[819] + MEM[92];
assign MEM[1214] = MEM[821] + MEM[557];
assign MEM[1215] = MEM[823] + MEM[30];
assign MEM[1216] = MEM[824] + MEM[4];
assign MEM[1217] = MEM[826] + MEM[319];
assign MEM[1218] = MEM[829] + MEM[679];
assign MEM[1219] = MEM[831] + MEM[726];
assign MEM[1220] = MEM[834] + MEM[274];
assign MEM[1221] = MEM[836] + MEM[801];
assign MEM[1222] = MEM[837] + MEM[251];
assign MEM[1223] = MEM[844] + MEM[451];
assign MEM[1224] = MEM[854] + MEM[366];
assign MEM[1225] = MEM[873] + MEM[589];
assign MEM[1226] = MEM[907] + MEM[717];
assign MEM[1227] = MEM[915] + MEM[650];
assign MEM[1228] = MEM[36] + MEM[763];
assign MEM[1229] = MEM[53] + MEM[742];
assign MEM[1230] = MEM[56] + MEM[699];
assign MEM[1231] = MEM[67] + MEM[852];
assign MEM[1232] = MEM[72] + MEM[527];
assign MEM[1233] = MEM[78] + MEM[603];
assign MEM[1234] = MEM[90] + MEM[147];
assign MEM[1235] = MEM[91] + MEM[745];
assign MEM[1236] = MEM[98] + MEM[294];
assign MEM[1237] = MEM[109] + MEM[746];
assign MEM[1238] = MEM[113] + MEM[157];
assign MEM[1239] = MEM[114] + MEM[695];
assign MEM[1240] = MEM[115] + MEM[220];
assign MEM[1241] = MEM[138] + MEM[803];
assign MEM[1242] = MEM[140] + MEM[792];
assign MEM[1243] = MEM[144] + MEM[527];
assign MEM[1244] = MEM[145] + MEM[144];
assign MEM[1245] = MEM[151] + MEM[849];
assign MEM[1246] = MEM[154] + MEM[641];
assign MEM[1247] = MEM[160] + MEM[229];
assign MEM[1248] = MEM[176] + MEM[493];
assign MEM[1249] = MEM[177] + MEM[530];
assign MEM[1250] = MEM[181] + MEM[355];
assign MEM[1251] = MEM[188] + MEM[146];
assign MEM[1252] = MEM[204] + MEM[551];
assign MEM[1253] = MEM[214] + MEM[870];
assign MEM[1254] = MEM[219] + MEM[625];
assign MEM[1255] = MEM[221] + MEM[567];
assign MEM[1256] = MEM[222] + MEM[662];
assign MEM[1257] = MEM[237] + MEM[261];
assign MEM[1258] = MEM[253] + MEM[519];
assign MEM[1259] = MEM[260] + MEM[771];
assign MEM[1260] = MEM[263] + MEM[203];
assign MEM[1261] = MEM[267] + MEM[73];
assign MEM[1262] = MEM[268] + MEM[514];
assign MEM[1263] = MEM[295] + MEM[777];
assign MEM[1264] = MEM[302] + MEM[733];
assign MEM[1265] = MEM[304] + MEM[866];
assign MEM[1266] = MEM[306] + MEM[182];
assign MEM[1267] = MEM[307] + MEM[710];
assign MEM[1268] = MEM[309] + MEM[340];
assign MEM[1269] = MEM[327] + MEM[464];
assign MEM[1270] = MEM[331] + MEM[460];
assign MEM[1271] = MEM[342] + MEM[428];
assign MEM[1272] = MEM[350] + MEM[523];
assign MEM[1273] = MEM[363] + MEM[667];
assign MEM[1274] = MEM[367] + MEM[43];
assign MEM[1275] = MEM[370] + MEM[855];
assign MEM[1276] = MEM[373] + MEM[660];
assign MEM[1277] = MEM[379] + MEM[814];
assign MEM[1278] = MEM[387] + MEM[684];
assign MEM[1279] = MEM[396] + MEM[458];
assign MEM[1280] = MEM[399] + MEM[672];
assign MEM[1281] = MEM[403] + MEM[841];
assign MEM[1282] = MEM[415] + MEM[754];
assign MEM[1283] = MEM[430] + MEM[29];
assign MEM[1284] = MEM[447] + MEM[532];
assign MEM[1285] = MEM[452] + MEM[1041];
assign MEM[1286] = MEM[459] + MEM[838];
assign MEM[1287] = MEM[463] + MEM[623];
assign MEM[1288] = MEM[465] + MEM[508];
assign MEM[1289] = MEM[480] + MEM[718];
assign MEM[1290] = MEM[487] + MEM[622];
assign MEM[1291] = MEM[501] + MEM[531];
assign MEM[1292] = MEM[503] + MEM[822];
assign MEM[1293] = MEM[523] + MEM[848];
assign MEM[1294] = MEM[526] + MEM[664];
assign MEM[1295] = MEM[528] + MEM[753];
assign MEM[1296] = MEM[535] + MEM[762];
assign MEM[1297] = MEM[538] + MEM[175];
assign MEM[1298] = MEM[548] + MEM[673];
assign MEM[1299] = MEM[550] + MEM[138];
assign MEM[1300] = MEM[550] + MEM[820];
assign MEM[1301] = MEM[558] + MEM[732];
assign MEM[1302] = MEM[562] + MEM[748];
assign MEM[1303] = MEM[579] + MEM[712];
assign MEM[1304] = MEM[582] + MEM[843];
assign MEM[1305] = MEM[588] + MEM[577];
assign MEM[1306] = MEM[591] + MEM[856];
assign MEM[1307] = MEM[599] + MEM[325];
assign MEM[1308] = MEM[601] + MEM[808];
assign MEM[1309] = MEM[612] + MEM[616];
assign MEM[1310] = MEM[615] + MEM[696];
assign MEM[1311] = MEM[630] + MEM[703];
assign MEM[1312] = MEM[635] + MEM[734];
assign MEM[1313] = MEM[640] + MEM[163];
assign MEM[1314] = MEM[643] + MEM[858];
assign MEM[1315] = MEM[644] + MEM[833];
assign MEM[1316] = MEM[653] + MEM[775];
assign MEM[1317] = MEM[654] + MEM[697];
assign MEM[1318] = MEM[655] + MEM[702];
assign MEM[1319] = MEM[659] + MEM[61];
assign MEM[1320] = MEM[667] + MEM[674];
assign MEM[1321] = MEM[675] + MEM[718];
assign MEM[1322] = MEM[677] + MEM[111];
assign MEM[1323] = MEM[689] + MEM[517];
assign MEM[1324] = MEM[711] + MEM[303];
assign MEM[1325] = MEM[715] + MEM[781];
assign MEM[1326] = MEM[716] + MEM[760];
assign MEM[1327] = MEM[720] + MEM[774];
assign MEM[1328] = MEM[723] + MEM[757];
assign MEM[1329] = MEM[730] + MEM[651];
assign MEM[1330] = MEM[738] + MEM[703];
assign MEM[1331] = MEM[741] + MEM[236];
assign MEM[1332] = MEM[743] + MEM[818];
assign MEM[1333] = MEM[748] + MEM[683];
assign MEM[1334] = MEM[749] + MEM[124];
assign MEM[1335] = MEM[750] + MEM[821];
assign MEM[1336] = MEM[751] + MEM[808];
assign MEM[1337] = MEM[754] + MEM[241];
assign MEM[1338] = MEM[755] + MEM[776];
assign MEM[1339] = MEM[758] + MEM[42];
assign MEM[1340] = MEM[759] + MEM[521];
assign MEM[1341] = MEM[764] + MEM[116];
assign MEM[1342] = MEM[766] + MEM[839];
assign MEM[1343] = MEM[769] + MEM[817];
assign MEM[1344] = MEM[770] + MEM[507];
assign MEM[1345] = MEM[779] + MEM[841];
assign MEM[1346] = MEM[780] + MEM[483];
assign MEM[1347] = MEM[782] + MEM[641];
assign MEM[1348] = MEM[786] + MEM[115];
assign MEM[1349] = MEM[787] + MEM[197];
assign MEM[1350] = MEM[790] + MEM[888];
assign MEM[1351] = MEM[797] + MEM[832];
assign MEM[1352] = MEM[800] + MEM[861];
assign MEM[1353] = MEM[805] + MEM[912];
assign MEM[1354] = MEM[810] + MEM[93];
assign MEM[1355] = MEM[832] + MEM[785];
assign MEM[1356] = MEM[840] + MEM[330];
assign MEM[1357] = MEM[842] + MEM[597];
assign MEM[1358] = MEM[845] + MEM[761];
assign MEM[1359] = MEM[850] + MEM[867];
assign MEM[1360] = MEM[851] + MEM[798];
assign MEM[1361] = MEM[857] + MEM[247];
assign MEM[1362] = MEM[859] + MEM[890];
assign MEM[1363] = MEM[860] + MEM[45];
assign MEM[1364] = MEM[862] + MEM[239];
assign MEM[1365] = MEM[868] + MEM[332];
assign MEM[1366] = MEM[872] + MEM[766];
assign MEM[1367] = MEM[874] + MEM[486];
assign MEM[1368] = MEM[879] + MEM[374];
assign MEM[1369] = MEM[882] + MEM[791];
assign MEM[1370] = MEM[885] + MEM[506];
assign MEM[1371] = MEM[908] + MEM[709];
assign MEM[1372] = MEM[948] + MEM[984];
assign MEM[1373] = MEM[1233] + MEM[604];
assign MEM[1374] = MEM[1259] + MEM[987];
assign MEM[1375] = MEM[1275] + MEM[1130];
assign MEM[1376] = MEM[2] + MEM[589];
assign MEM[1377] = MEM[3] + MEM[125];
assign MEM[1378] = MEM[4] + MEM[770];
assign MEM[1379] = MEM[5] + MEM[101];
assign MEM[1380] = MEM[7] + MEM[477];
assign MEM[1381] = MEM[10] + MEM[783];
assign MEM[1382] = MEM[11] + MEM[501];
assign MEM[1383] = MEM[12] + MEM[64];
assign MEM[1384] = MEM[13] + MEM[599];
assign MEM[1385] = MEM[18] + MEM[83];
assign MEM[1386] = MEM[19] + MEM[638];
assign MEM[1387] = MEM[21] + MEM[157];
assign MEM[1388] = MEM[26] + MEM[218];
assign MEM[1389] = MEM[27] + MEM[460];
assign MEM[1390] = MEM[31] + MEM[59];
assign MEM[1391] = MEM[34] + MEM[37];
assign MEM[1392] = MEM[35] + MEM[245];
assign MEM[1393] = MEM[36] + MEM[824];
assign MEM[1394] = MEM[38] + MEM[537];
assign MEM[1395] = MEM[39] + MEM[568];
assign MEM[1396] = MEM[44] + MEM[141];
assign MEM[1397] = MEM[47] + MEM[611];
assign MEM[1398] = MEM[50] + MEM[242];
assign MEM[1399] = MEM[53] + MEM[323];
assign MEM[1400] = MEM[56] + MEM[372];
assign MEM[1401] = MEM[57] + MEM[445];
assign MEM[1402] = MEM[58] + MEM[853];
assign MEM[1403] = MEM[60] + MEM[900];
assign MEM[1404] = MEM[62] + MEM[1048];
assign MEM[1405] = MEM[63] + MEM[178];
assign MEM[1406] = MEM[63] + MEM[930];
assign MEM[1407] = MEM[64] + MEM[654];
assign MEM[1408] = MEM[65] + MEM[617];
assign MEM[1409] = MEM[66] + MEM[272];
assign MEM[1410] = MEM[69] + MEM[191];
assign MEM[1411] = MEM[70] + MEM[889];
assign MEM[1412] = MEM[72] + MEM[288];
assign MEM[1413] = MEM[74] + MEM[450];
assign MEM[1414] = MEM[75] + MEM[348];
assign MEM[1415] = MEM[76] + MEM[364];
assign MEM[1416] = MEM[79] + MEM[474];
assign MEM[1417] = MEM[84] + MEM[939];
assign MEM[1418] = MEM[85] + MEM[386];
assign MEM[1419] = MEM[86] + MEM[278];
assign MEM[1420] = MEM[86] + MEM[575];
assign MEM[1421] = MEM[87] + MEM[277];
assign MEM[1422] = MEM[95] + MEM[762];
assign MEM[1423] = MEM[99] + MEM[570];
assign MEM[1424] = MEM[100] + MEM[590];
assign MEM[1425] = MEM[106] + MEM[291];
assign MEM[1426] = MEM[107] + MEM[757];
assign MEM[1427] = MEM[108] + MEM[165];
assign MEM[1428] = MEM[112] + MEM[275];
assign MEM[1429] = MEM[113] + MEM[979];
assign MEM[1430] = MEM[117] + MEM[143];
assign MEM[1431] = MEM[118] + MEM[179];
assign MEM[1432] = MEM[119] + MEM[669];
assign MEM[1433] = MEM[119] + MEM[1108];
assign MEM[1434] = MEM[122] + MEM[341];
assign MEM[1435] = MEM[123] + MEM[730];
assign MEM[1436] = MEM[130] + MEM[653];
assign MEM[1437] = MEM[131] + MEM[833];
assign MEM[1438] = MEM[132] + MEM[149];
assign MEM[1439] = MEM[133] + MEM[563];
assign MEM[1440] = MEM[134] + MEM[287];
assign MEM[1441] = MEM[141] + MEM[744];
assign MEM[1442] = MEM[145] + MEM[884];
assign MEM[1443] = MEM[155] + MEM[839];
assign MEM[1444] = MEM[156] + MEM[418];
assign MEM[1445] = MEM[158] + MEM[307];
assign MEM[1446] = MEM[161] + MEM[799];
assign MEM[1447] = MEM[162] + MEM[298];
assign MEM[1448] = MEM[167] + MEM[495];
assign MEM[1449] = MEM[171] + MEM[585];
assign MEM[1450] = MEM[173] + MEM[543];
assign MEM[1451] = MEM[174] + MEM[886];
assign MEM[1452] = MEM[176] + MEM[554];
assign MEM[1453] = MEM[178] + MEM[479];
assign MEM[1454] = MEM[180] + MEM[516];
assign MEM[1455] = MEM[181] + MEM[308];
assign MEM[1456] = MEM[185] + MEM[426];
assign MEM[1457] = MEM[186] + MEM[252];
assign MEM[1458] = MEM[187] + MEM[250];
assign MEM[1459] = MEM[189] + MEM[756];
assign MEM[1460] = MEM[190] + MEM[595];
assign MEM[1461] = MEM[194] + MEM[560];
assign MEM[1462] = MEM[195] + MEM[207];
assign MEM[1463] = MEM[196] + MEM[310];
assign MEM[1464] = MEM[199] + MEM[431];
assign MEM[1465] = MEM[201] + MEM[863];
assign MEM[1466] = MEM[202] + MEM[251];
assign MEM[1467] = MEM[204] + MEM[610];
assign MEM[1468] = MEM[206] + MEM[956];
assign MEM[1469] = MEM[210] + MEM[1190];
assign MEM[1470] = MEM[212] + MEM[365];
assign MEM[1471] = MEM[213] + MEM[622];
assign MEM[1472] = MEM[215] + MEM[476];
assign MEM[1473] = MEM[218] + MEM[1111];
assign MEM[1474] = MEM[219] + MEM[416];
assign MEM[1475] = MEM[222] + MEM[807];
assign MEM[1476] = MEM[223] + MEM[895];
assign MEM[1477] = MEM[227] + MEM[404];
assign MEM[1478] = MEM[228] + MEM[551];
assign MEM[1479] = MEM[230] + MEM[302];
assign MEM[1480] = MEM[231] + MEM[469];
assign MEM[1481] = MEM[233] + MEM[794];
assign MEM[1482] = MEM[234] + MEM[772];
assign MEM[1483] = MEM[235] + MEM[661];
assign MEM[1484] = MEM[238] + MEM[357];
assign MEM[1485] = MEM[238] + MEM[566];
assign MEM[1486] = MEM[240] + MEM[898];
assign MEM[1487] = MEM[242] + MEM[893];
assign MEM[1488] = MEM[243] + MEM[478];
assign MEM[1489] = MEM[245] + MEM[727];
assign MEM[1490] = MEM[246] + MEM[649];
assign MEM[1491] = MEM[253] + MEM[938];
assign MEM[1492] = MEM[254] + MEM[586];
assign MEM[1493] = MEM[259] + MEM[467];
assign MEM[1494] = MEM[262] + MEM[746];
assign MEM[1495] = MEM[266] + MEM[814];
assign MEM[1496] = MEM[267] + MEM[864];
assign MEM[1497] = MEM[269] + MEM[847];
assign MEM[1498] = MEM[273] + MEM[1029];
assign MEM[1499] = MEM[274] + MEM[951];
assign MEM[1500] = MEM[279] + MEM[371];
assign MEM[1501] = MEM[283] + MEM[397];
assign MEM[1502] = MEM[284] + MEM[962];
assign MEM[1503] = MEM[286] + MEM[333];
assign MEM[1504] = MEM[288] + MEM[289];
assign MEM[1505] = MEM[290] + MEM[779];
assign MEM[1506] = MEM[292] + MEM[851];
assign MEM[1507] = MEM[293] + MEM[414];
assign MEM[1508] = MEM[296] + MEM[546];
assign MEM[1509] = MEM[298] + MEM[865];
assign MEM[1510] = MEM[301] + MEM[389];
assign MEM[1511] = MEM[301] + MEM[929];
assign MEM[1512] = MEM[305] + MEM[608];
assign MEM[1513] = MEM[314] + MEM[338];
assign MEM[1514] = MEM[315] + MEM[949];
assign MEM[1515] = MEM[318] + MEM[806];
assign MEM[1516] = MEM[322] + MEM[406];
assign MEM[1517] = MEM[324] + MEM[986];
assign MEM[1518] = MEM[326] + MEM[343];
assign MEM[1519] = MEM[331] + MEM[796];
assign MEM[1520] = MEM[334] + MEM[871];
assign MEM[1521] = MEM[334] + MEM[1139];
assign MEM[1522] = MEM[335] + MEM[883];
assign MEM[1523] = MEM[336] + MEM[806];
assign MEM[1524] = MEM[339] + MEM[765];
assign MEM[1525] = MEM[340] + MEM[244];
assign MEM[1526] = MEM[346] + MEM[765];
assign MEM[1527] = MEM[346] + MEM[785];
assign MEM[1528] = MEM[349] + MEM[390];
assign MEM[1529] = MEM[350] + MEM[571];
assign MEM[1530] = MEM[351] + MEM[88];
assign MEM[1531] = MEM[354] + MEM[696];
assign MEM[1532] = MEM[355] + MEM[584];
assign MEM[1533] = MEM[358] + MEM[576];
assign MEM[1534] = MEM[359] + MEM[633];
assign MEM[1535] = MEM[367] + MEM[436];
assign MEM[1536] = MEM[367] + MEM[695];
assign MEM[1537] = MEM[375] + MEM[545];
assign MEM[1538] = MEM[378] + MEM[788];
assign MEM[1539] = MEM[382] + MEM[402];
assign MEM[1540] = MEM[388] + MEM[559];
assign MEM[1541] = MEM[391] + MEM[544];
assign MEM[1542] = MEM[394] + MEM[699];
assign MEM[1543] = MEM[394] + MEM[891];
assign MEM[1544] = MEM[404] + MEM[997];
assign MEM[1545] = MEM[405] + MEM[587];
assign MEM[1546] = MEM[407] + MEM[540];
assign MEM[1547] = MEM[407] + MEM[1255];
assign MEM[1548] = MEM[418] + MEM[1044];
assign MEM[1549] = MEM[420] + MEM[773];
assign MEM[1550] = MEM[427] + MEM[583];
assign MEM[1551] = MEM[428] + MEM[659];
assign MEM[1552] = MEM[435] + MEM[728];
assign MEM[1553] = MEM[437] + MEM[549];
assign MEM[1554] = MEM[439] + MEM[792];
assign MEM[1555] = MEM[440] + MEM[655];
assign MEM[1556] = MEM[443] + MEM[582];
assign MEM[1557] = MEM[446] + MEM[818];
assign MEM[1558] = MEM[446] + MEM[933];
assign MEM[1559] = MEM[448] + MEM[485];
assign MEM[1560] = MEM[449] + MEM[475];
assign MEM[1561] = MEM[450] + MEM[917];
assign MEM[1562] = MEM[451] + MEM[455];
assign MEM[1563] = MEM[453] + MEM[772];
assign MEM[1564] = MEM[454] + MEM[618];
assign MEM[1565] = MEM[457] + MEM[592];
assign MEM[1566] = MEM[458] + MEM[676];
assign MEM[1567] = MEM[464] + MEM[819];
assign MEM[1568] = MEM[465] + MEM[564];
assign MEM[1569] = MEM[466] + MEM[658];
assign MEM[1570] = MEM[467] + MEM[1050];
assign MEM[1571] = MEM[468] + MEM[188];
assign MEM[1572] = MEM[468] + MEM[634];
assign MEM[1573] = MEM[469] + MEM[852];
assign MEM[1574] = MEM[470] + MEM[627];
assign MEM[1575] = MEM[477] + MEM[921];
assign MEM[1576] = MEM[479] + MEM[1166];
assign MEM[1577] = MEM[481] + MEM[585];
assign MEM[1578] = MEM[482] + MEM[35];
assign MEM[1579] = MEM[484] + MEM[660];
assign MEM[1580] = MEM[484] + MEM[676];
assign MEM[1581] = MEM[490] + MEM[628];
assign MEM[1582] = MEM[491] + MEM[886];
assign MEM[1583] = MEM[492] + MEM[154];
assign MEM[1584] = MEM[499] + MEM[1145];
assign MEM[1585] = MEM[500] + MEM[1097];
assign MEM[1586] = MEM[509] + MEM[894];
assign MEM[1587] = MEM[510] + MEM[1002];
assign MEM[1588] = MEM[511] + MEM[927];
assign MEM[1589] = MEM[518] + MEM[1039];
assign MEM[1590] = MEM[520] + MEM[877];
assign MEM[1591] = MEM[522] + MEM[816];
assign MEM[1592] = MEM[522] + MEM[947];
assign MEM[1593] = MEM[528] + MEM[1113];
assign MEM[1594] = MEM[529] + MEM[732];
assign MEM[1595] = MEM[530] + MEM[687];
assign MEM[1596] = MEM[531] + MEM[1035];
assign MEM[1597] = MEM[533] + MEM[838];
assign MEM[1598] = MEM[533] + MEM[950];
assign MEM[1599] = MEM[534] + MEM[410];
assign MEM[1600] = MEM[535] + MEM[946];
assign MEM[1601] = MEM[535] + MEM[983];
assign MEM[1602] = MEM[537] + MEM[828];
assign MEM[1603] = MEM[539] + MEM[720];
assign MEM[1604] = MEM[542] + MEM[804];
assign MEM[1605] = MEM[543] + MEM[670];
assign MEM[1606] = MEM[551] + MEM[782];
assign MEM[1607] = MEM[553] + MEM[925];
assign MEM[1608] = MEM[554] + MEM[673];
assign MEM[1609] = MEM[555] + MEM[624];
assign MEM[1610] = MEM[556] + MEM[691];
assign MEM[1611] = MEM[557] + MEM[867];
assign MEM[1612] = MEM[563] + MEM[863];
assign MEM[1613] = MEM[565] + MEM[822];
assign MEM[1614] = MEM[574] + MEM[365];
assign MEM[1615] = MEM[576] + MEM[705];
assign MEM[1616] = MEM[580] + MEM[922];
assign MEM[1617] = MEM[581] + MEM[737];
assign MEM[1618] = MEM[586] + MEM[876];
assign MEM[1619] = MEM[594] + MEM[906];
assign MEM[1620] = MEM[600] + MEM[1077];
assign MEM[1621] = MEM[602] + MEM[429];
assign MEM[1622] = MEM[605] + MEM[789];
assign MEM[1623] = MEM[606] + MEM[613];
assign MEM[1624] = MEM[607] + MEM[833];
assign MEM[1625] = MEM[612] + MEM[985];
assign MEM[1626] = MEM[614] + MEM[977];
assign MEM[1627] = MEM[614] + MEM[1092];
assign MEM[1628] = MEM[619] + MEM[715];
assign MEM[1629] = MEM[620] + MEM[771];
assign MEM[1630] = MEM[621] + MEM[1045];
assign MEM[1631] = MEM[623] + MEM[802];
assign MEM[1632] = MEM[625] + MEM[939];
assign MEM[1633] = MEM[635] + MEM[1065];
assign MEM[1634] = MEM[636] + MEM[883];
assign MEM[1635] = MEM[636] + MEM[896];
assign MEM[1636] = MEM[639] + MEM[827];
assign MEM[1637] = MEM[642] + MEM[913];
assign MEM[1638] = MEM[642] + MEM[1122];
assign MEM[1639] = MEM[645] + MEM[918];
assign MEM[1640] = MEM[646] + MEM[856];
assign MEM[1641] = MEM[650] + MEM[710];
assign MEM[1642] = MEM[655] + MEM[717];
assign MEM[1643] = MEM[664] + MEM[707];
assign MEM[1644] = MEM[665] + MEM[778];
assign MEM[1645] = MEM[666] + MEM[682];
assign MEM[1646] = MEM[667] + MEM[686];
assign MEM[1647] = MEM[668] + MEM[850];
assign MEM[1648] = MEM[669] + MEM[1006];
assign MEM[1649] = MEM[675] + MEM[836];
assign MEM[1650] = MEM[677] + MEM[648];
assign MEM[1651] = MEM[677] + MEM[866];
assign MEM[1652] = MEM[682] + MEM[813];
assign MEM[1653] = MEM[684] + MEM[880];
assign MEM[1654] = MEM[685] + MEM[1180];
assign MEM[1655] = MEM[687] + MEM[842];
assign MEM[1656] = MEM[689] + MEM[413];
assign MEM[1657] = MEM[692] + MEM[889];
assign MEM[1658] = MEM[692] + MEM[903];
assign MEM[1659] = MEM[700] + MEM[835];
assign MEM[1660] = MEM[701] + MEM[952];
assign MEM[1661] = MEM[704] + MEM[271];
assign MEM[1662] = MEM[708] + MEM[762];
assign MEM[1663] = MEM[714] + MEM[444];
assign MEM[1664] = MEM[716] + MEM[937];
assign MEM[1665] = MEM[719] + MEM[783];
assign MEM[1666] = MEM[723] + MEM[793];
assign MEM[1667] = MEM[725] + MEM[1568];
assign MEM[1668] = MEM[726] + MEM[861];
assign MEM[1669] = MEM[729] + MEM[909];
assign MEM[1670] = MEM[733] + MEM[999];
assign MEM[1671] = MEM[733] + MEM[1220];
assign MEM[1672] = MEM[734] + MEM[795];
assign MEM[1673] = MEM[739] + MEM[853];
assign MEM[1674] = MEM[741] + MEM[875];
assign MEM[1675] = MEM[742] + MEM[481];
assign MEM[1676] = MEM[745] + MEM[874];
assign MEM[1677] = MEM[749] + MEM[826];
assign MEM[1678] = MEM[753] + MEM[610];
assign MEM[1679] = MEM[755] + MEM[799];
assign MEM[1680] = MEM[758] + MEM[1049];
assign MEM[1681] = MEM[759] + MEM[1090];
assign MEM[1682] = MEM[763] + MEM[944];
assign MEM[1683] = MEM[768] + MEM[981];
assign MEM[1684] = MEM[769] + MEM[1042];
assign MEM[1685] = MEM[773] + MEM[901];
assign MEM[1686] = MEM[781] + MEM[980];
assign MEM[1687] = MEM[786] + MEM[843];
assign MEM[1688] = MEM[791] + MEM[967];
assign MEM[1689] = MEM[793] + MEM[869];
assign MEM[1690] = MEM[794] + MEM[973];
assign MEM[1691] = MEM[807] + MEM[936];
assign MEM[1692] = MEM[809] + MEM[1031];
assign MEM[1693] = MEM[810] + MEM[904];
assign MEM[1694] = MEM[810] + MEM[1056];
assign MEM[1695] = MEM[811] + MEM[812];
assign MEM[1696] = MEM[811] + MEM[1051];
assign MEM[1697] = MEM[815] + MEM[842];
assign MEM[1698] = MEM[818] + MEM[971];
assign MEM[1699] = MEM[823] + MEM[200];
assign MEM[1700] = MEM[825] + MEM[937];
assign MEM[1701] = MEM[826] + MEM[1138];
assign MEM[1702] = MEM[829] + MEM[15];
assign MEM[1703] = MEM[830] + MEM[1021];
assign MEM[1704] = MEM[837] + MEM[1046];
assign MEM[1705] = MEM[844] + MEM[921];
assign MEM[1706] = MEM[846] + MEM[902];
assign MEM[1707] = MEM[847] + MEM[949];
assign MEM[1708] = MEM[848] + MEM[1116];
assign MEM[1709] = MEM[852] + MEM[878];
assign MEM[1710] = MEM[854] + MEM[640];
assign MEM[1711] = MEM[855] + MEM[975];
assign MEM[1712] = MEM[860] + MEM[815];
assign MEM[1713] = MEM[864] + MEM[942];
assign MEM[1714] = MEM[869] + MEM[887];
assign MEM[1715] = MEM[871] + MEM[911];
assign MEM[1716] = MEM[875] + MEM[1124];
assign MEM[1717] = MEM[876] + MEM[1000];
assign MEM[1718] = MEM[880] + MEM[932];
assign MEM[1719] = MEM[881] + MEM[1025];
assign MEM[1720] = MEM[890] + MEM[542];
assign MEM[1721] = MEM[892] + MEM[637];
assign MEM[1722] = MEM[894] + MEM[1093];
assign MEM[1723] = MEM[897] + MEM[968];
assign MEM[1724] = MEM[905] + MEM[923];
assign MEM[1725] = MEM[910] + MEM[738];
assign MEM[1726] = MEM[911] + MEM[951];
assign MEM[1727] = MEM[914] + MEM[964];
assign MEM[1728] = MEM[916] + MEM[1198];
assign MEM[1729] = MEM[919] + MEM[172];
assign MEM[1730] = MEM[919] + MEM[1007];
assign MEM[1731] = MEM[920] + MEM[434];
assign MEM[1732] = MEM[924] + MEM[927];
assign MEM[1733] = MEM[926] + MEM[972];
assign MEM[1734] = MEM[928] + MEM[1036];
assign MEM[1735] = MEM[931] + MEM[969];
assign MEM[1736] = MEM[932] + MEM[933];
assign MEM[1737] = MEM[934] + MEM[978];
assign MEM[1738] = MEM[935] + MEM[1022];
assign MEM[1739] = MEM[940] + MEM[1132];
assign MEM[1740] = MEM[941] + MEM[1071];
assign MEM[1741] = MEM[943] + MEM[1073];
assign MEM[1742] = MEM[945] + MEM[804];
assign MEM[1743] = MEM[953] + MEM[1009];
assign MEM[1744] = MEM[954] + MEM[1070];
assign MEM[1745] = MEM[960] + MEM[905];
assign MEM[1746] = MEM[963] + MEM[712];
assign MEM[1747] = MEM[966] + MEM[545];
assign MEM[1748] = MEM[970] + MEM[1063];
assign MEM[1749] = MEM[970] + MEM[1064];
assign MEM[1750] = MEM[972] + MEM[1224];
assign MEM[1751] = MEM[976] + MEM[926];
assign MEM[1752] = MEM[988] + MEM[1151];
assign MEM[1753] = MEM[990] + MEM[849];
assign MEM[1754] = MEM[991] + MEM[1019];
assign MEM[1755] = MEM[991] + MEM[1150];
assign MEM[1756] = MEM[994] + MEM[891];
assign MEM[1757] = MEM[995] + MEM[423];
assign MEM[1758] = MEM[996] + MEM[629];
assign MEM[1759] = MEM[998] + MEM[1013];
assign MEM[1760] = MEM[1001] + MEM[750];
assign MEM[1761] = MEM[1002] + MEM[1174];
assign MEM[1762] = MEM[1003] + MEM[1112];
assign MEM[1763] = MEM[1006] + MEM[1160];
assign MEM[1764] = MEM[1010] + MEM[1176];
assign MEM[1765] = MEM[1010] + MEM[1733];
assign MEM[1766] = MEM[1011] + MEM[702];
assign MEM[1767] = MEM[1014] + MEM[892];
assign MEM[1768] = MEM[1014] + MEM[1033];
assign MEM[1769] = MEM[1015] + MEM[1047];
assign MEM[1770] = MEM[1024] + MEM[347];
assign MEM[1771] = MEM[1029] + MEM[1168];
assign MEM[1772] = MEM[1032] + MEM[1037];
assign MEM[1773] = MEM[1040] + MEM[1131];
assign MEM[1774] = MEM[1043] + MEM[1194];
assign MEM[1775] = MEM[1053] + MEM[1159];
assign MEM[1776] = MEM[1054] + MEM[732];
assign MEM[1777] = MEM[1059] + MEM[857];
assign MEM[1778] = MEM[1060] + MEM[1203];
assign MEM[1779] = MEM[1061] + MEM[1016];
assign MEM[1780] = MEM[1064] + MEM[1038];
assign MEM[1781] = MEM[1067] + MEM[1055];
assign MEM[1782] = MEM[1068] + MEM[1078];
assign MEM[1783] = MEM[1076] + MEM[1104];
assign MEM[1784] = MEM[1086] + MEM[822];
assign MEM[1785] = MEM[1105] + MEM[1084];
assign MEM[1786] = MEM[1128] + MEM[882];
assign MEM[1787] = MEM[1140] + MEM[1125];
assign MEM[1788] = MEM[1142] + MEM[929];
assign MEM[1789] = MEM[1149] + MEM[961];
assign MEM[1790] = MEM[1155] + MEM[862];
assign MEM[1791] = MEM[1161] + MEM[150];
assign MEM[1792] = MEM[1164] + MEM[965];
assign MEM[1793] = MEM[1171] + MEM[1178];
assign MEM[1794] = MEM[1191] + MEM[1156];
assign MEM[1795] = MEM[1193] + MEM[938];
assign MEM[1796] = MEM[1221] + MEM[1034];
assign MEM[1797] = MEM[1226] + MEM[884];
assign MEM[1798] = MEM[1227] + MEM[1153];
assign MEM[1799] = MEM[1230] + MEM[840];
assign MEM[1800] = MEM[1237] + MEM[1057];
assign MEM[1801] = MEM[1298] + MEM[351];
assign MEM[1802] = MEM[1300] + MEM[922];
assign MEM[1803] = MEM[1386] + MEM[1107];
assign MEM[1804] = MEM[1417] + MEM[1114];
assign MEM[1805] = MEM[1420] + MEM[1026];
assign MEM[1806] = MEM[1462] + MEM[1664];
assign MEM[1807] = MEM[1466] + MEM[1075];
assign MEM[1808] = MEM[1501] + MEM[878];
assign MEM[1809] = MEM[1503] + MEM[1136];
assign MEM[1810] = MEM[1559] + MEM[1087];
assign MEM[1811] = MEM[1625] + MEM[1117];
assign MEM[1812] = MEM[1639] + MEM[1768];
assign MEM[1813] = MEM[1680] + MEM[1201];
assign MEM[1814] = MEM[1686] + MEM[1005];
assign MEM[1815] = MEM[1736] + MEM[992];
assign MEM[1816] = MEM[2] + MEM[1373];
assign MEM[1817] = MEM[3] + MEM[163];
assign MEM[1818] = MEM[6] + MEM[73];
assign MEM[1819] = MEM[6] + MEM[579];
assign MEM[1820] = MEM[7] + MEM[668];
assign MEM[1821] = MEM[11] + MEM[899];
assign MEM[1822] = MEM[12] + MEM[508];
assign MEM[1823] = MEM[13] + MEM[606];
assign MEM[1824] = MEM[14] + MEM[801];
assign MEM[1825] = MEM[14] + MEM[1213];
assign MEM[1826] = MEM[15] + MEM[946];
assign MEM[1827] = MEM[17] + MEM[1081];
assign MEM[1828] = MEM[18] + MEM[427];
assign MEM[1829] = MEM[19] + MEM[221];
assign MEM[1830] = MEM[20] + MEM[308];
assign MEM[1831] = MEM[20] + MEM[324];
assign MEM[1832] = MEM[21] + MEM[993];
assign MEM[1833] = MEM[22] + MEM[306];
assign MEM[1834] = MEM[23] + MEM[893];
assign MEM[1835] = MEM[26] + MEM[90];
assign MEM[1836] = MEM[28] + MEM[233];
assign MEM[1837] = MEM[28] + MEM[802];
assign MEM[1838] = MEM[29] + MEM[71];
assign MEM[1839] = MEM[31] + MEM[564];
assign MEM[1840] = MEM[34] + MEM[656];
assign MEM[1841] = MEM[36] + MEM[727];
assign MEM[1842] = MEM[37] + MEM[48];
assign MEM[1843] = MEM[38] + MEM[626];
assign MEM[1844] = MEM[43] + MEM[441];
assign MEM[1845] = MEM[44] + MEM[887];
assign MEM[1846] = MEM[45] + MEM[930];
assign MEM[1847] = MEM[46] + MEM[57];
assign MEM[1848] = MEM[47] + MEM[1123];
assign MEM[1849] = MEM[50] + MEM[777];
assign MEM[1850] = MEM[51] + MEM[110];
assign MEM[1851] = MEM[51] + MEM[1098];
assign MEM[1852] = MEM[52] + MEM[158];
assign MEM[1853] = MEM[52] + MEM[430];
assign MEM[1854] = MEM[53] + MEM[1711];
assign MEM[1855] = MEM[55] + MEM[568];
assign MEM[1856] = MEM[58] + MEM[630];
assign MEM[1857] = MEM[59] + MEM[328];
assign MEM[1858] = MEM[59] + MEM[868];
assign MEM[1859] = MEM[60] + MEM[94];
assign MEM[1860] = MEM[61] + MEM[955];
assign MEM[1861] = MEM[62] + MEM[419];
assign MEM[1862] = MEM[64] + MEM[729];
assign MEM[1863] = MEM[66] + MEM[259];
assign MEM[1864] = MEM[66] + MEM[713];
assign MEM[1865] = MEM[67] + MEM[944];
assign MEM[1866] = MEM[68] + MEM[1042];
assign MEM[1867] = MEM[69] + MEM[688];
assign MEM[1868] = MEM[70] + MEM[931];
assign MEM[1869] = MEM[71] + MEM[963];
assign MEM[1870] = MEM[72] + MEM[1185];
assign MEM[1871] = MEM[75] + MEM[373];
assign MEM[1872] = MEM[77] + MEM[380];
assign MEM[1873] = MEM[77] + MEM[957];
assign MEM[1874] = MEM[78] + MEM[555];
assign MEM[1875] = MEM[79] + MEM[463];
assign MEM[1876] = MEM[82] + MEM[103];
assign MEM[1877] = MEM[83] + MEM[788];
assign MEM[1878] = MEM[85] + MEM[1151];
assign MEM[1879] = MEM[87] + MEM[1023];
assign MEM[1880] = MEM[88] + MEM[1535];
assign MEM[1881] = MEM[89] + MEM[452];
assign MEM[1882] = MEM[89] + MEM[1094];
assign MEM[1883] = MEM[90] + MEM[312];
assign MEM[1884] = MEM[90] + MEM[775];
assign MEM[1885] = MEM[93] + MEM[1239];
assign MEM[1886] = MEM[94] + MEM[461];
assign MEM[1887] = MEM[95] + MEM[398];
assign MEM[1888] = MEM[96] + MEM[778];
assign MEM[1889] = MEM[99] + MEM[1018];
assign MEM[1890] = MEM[101] + MEM[686];
assign MEM[1891] = MEM[102] + MEM[1106];
assign MEM[1892] = MEM[103] + MEM[1231];
assign MEM[1893] = MEM[106] + MEM[1121];
assign MEM[1894] = MEM[107] + MEM[753];
assign MEM[1895] = MEM[108] + MEM[803];
assign MEM[1896] = MEM[110] + MEM[880];
assign MEM[1897] = MEM[112] + MEM[400];
assign MEM[1898] = MEM[113] + MEM[945];
assign MEM[1899] = MEM[114] + MEM[877];
assign MEM[1900] = MEM[115] + MEM[1212];
assign MEM[1901] = MEM[117] + MEM[879];
assign MEM[1902] = MEM[117] + MEM[297];
assign MEM[1903] = MEM[118] + MEM[760];
assign MEM[1904] = MEM[118] + MEM[1182];
assign MEM[1905] = MEM[122] + MEM[1341];
assign MEM[1906] = MEM[123] + MEM[971];
assign MEM[1907] = MEM[124] + MEM[1152];
assign MEM[1908] = MEM[125] + MEM[1297];
assign MEM[1909] = MEM[126] + MEM[205];
assign MEM[1910] = MEM[127] + MEM[355];
assign MEM[1911] = MEM[130] + MEM[673];
assign MEM[1912] = MEM[131] + MEM[270];
assign MEM[1913] = MEM[132] + MEM[1078];
assign MEM[1914] = MEM[133] + MEM[1289];
assign MEM[1915] = MEM[134] + MEM[1729];
assign MEM[1916] = MEM[135] + MEM[295];
assign MEM[1917] = MEM[135] + MEM[375];
assign MEM[1918] = MEM[142] + MEM[166];
assign MEM[1919] = MEM[143] + MEM[390];
assign MEM[1920] = MEM[147] + MEM[641];
assign MEM[1921] = MEM[148] + MEM[199];
assign MEM[1922] = MEM[148] + MEM[438];
assign MEM[1923] = MEM[149] + MEM[383];
assign MEM[1924] = MEM[155] + MEM[923];
assign MEM[1925] = MEM[156] + MEM[1025];
assign MEM[1926] = MEM[157] + MEM[305];
assign MEM[1927] = MEM[159] + MEM[1367];
assign MEM[1928] = MEM[160] + MEM[1033];
assign MEM[1929] = MEM[161] + MEM[513];
assign MEM[1930] = MEM[162] + MEM[617];
assign MEM[1931] = MEM[165] + MEM[437];
assign MEM[1932] = MEM[167] + MEM[211];
assign MEM[1933] = MEM[173] + MEM[494];
assign MEM[1934] = MEM[176] + MEM[572];
assign MEM[1935] = MEM[177] + MEM[395];
assign MEM[1936] = MEM[180] + MEM[657];
assign MEM[1937] = MEM[181] + MEM[859];
assign MEM[1938] = MEM[182] + MEM[751];
assign MEM[1939] = MEM[183] + MEM[198];
assign MEM[1940] = MEM[183] + MEM[909];
assign MEM[1941] = MEM[185] + MEM[548];
assign MEM[1942] = MEM[186] + MEM[608];
assign MEM[1943] = MEM[187] + MEM[899];
assign MEM[1944] = MEM[190] + MEM[229];
assign MEM[1945] = MEM[191] + MEM[1254];
assign MEM[1946] = MEM[192] + MEM[1274];
assign MEM[1947] = MEM[195] + MEM[566];
assign MEM[1948] = MEM[196] + MEM[690];
assign MEM[1949] = MEM[197] + MEM[718];
assign MEM[1950] = MEM[198] + MEM[411];
assign MEM[1951] = MEM[201] + MEM[1008];
assign MEM[1952] = MEM[202] + MEM[414];
assign MEM[1953] = MEM[203] + MEM[260];
assign MEM[1954] = MEM[204] + MEM[553];
assign MEM[1955] = MEM[205] + MEM[1540];
assign MEM[1956] = MEM[206] + MEM[1009];
assign MEM[1957] = MEM[211] + MEM[671];
assign MEM[1958] = MEM[212] + MEM[402];
assign MEM[1959] = MEM[213] + MEM[1048];
assign MEM[1960] = MEM[214] + MEM[872];
assign MEM[1961] = MEM[215] + MEM[895];
assign MEM[1962] = MEM[217] + MEM[872];
assign MEM[1963] = MEM[219] + MEM[593];
assign MEM[1964] = MEM[220] + MEM[1256];
assign MEM[1965] = MEM[222] + MEM[712];
assign MEM[1966] = MEM[223] + MEM[1402];
assign MEM[1967] = MEM[227] + MEM[858];
assign MEM[1968] = MEM[228] + MEM[272];
assign MEM[1969] = MEM[229] + MEM[487];
assign MEM[1970] = MEM[231] + MEM[743];
assign MEM[1971] = MEM[232] + MEM[622];
assign MEM[1972] = MEM[234] + MEM[493];
assign MEM[1973] = MEM[235] + MEM[582];
assign MEM[1974] = MEM[236] + MEM[1096];
assign MEM[1975] = MEM[237] + MEM[1023];
assign MEM[1976] = MEM[239] + MEM[1290];
assign MEM[1977] = MEM[240] + MEM[790];
assign MEM[1978] = MEM[243] + MEM[442];
assign MEM[1979] = MEM[244] + MEM[420];
assign MEM[1980] = MEM[246] + MEM[888];
assign MEM[1981] = MEM[250] + MEM[293];
assign MEM[1982] = MEM[252] + MEM[1235];
assign MEM[1983] = MEM[255] + MEM[310];
assign MEM[1984] = MEM[255] + MEM[631];
assign MEM[1985] = MEM[258] + MEM[443];
assign MEM[1986] = MEM[261] + MEM[709];
assign MEM[1987] = MEM[262] + MEM[1101];
assign MEM[1988] = MEM[263] + MEM[1188];
assign MEM[1989] = MEM[266] + MEM[904];
assign MEM[1990] = MEM[268] + MEM[583];
assign MEM[1991] = MEM[270] + MEM[412];
assign MEM[1992] = MEM[275] + MEM[744];
assign MEM[1993] = MEM[276] + MEM[278];
assign MEM[1994] = MEM[277] + MEM[285];
assign MEM[1995] = MEM[278] + MEM[1037];
assign MEM[1996] = MEM[279] + MEM[1396];
assign MEM[1997] = MEM[283] + MEM[1128];
assign MEM[1998] = MEM[284] + MEM[1316];
assign MEM[1999] = MEM[286] + MEM[335];
assign MEM[2000] = MEM[287] + MEM[311];
assign MEM[2001] = MEM[289] + MEM[575];
assign MEM[2002] = MEM[291] + MEM[516];
assign MEM[2003] = MEM[292] + MEM[1144];
assign MEM[2004] = MEM[294] + MEM[774];
assign MEM[2005] = MEM[296] + MEM[601];
assign MEM[2006] = MEM[297] + MEM[326];
assign MEM[2007] = MEM[299] + MEM[657];
assign MEM[2008] = MEM[300] + MEM[1737];
assign MEM[2009] = MEM[302] + MEM[436];
assign MEM[2010] = MEM[303] + MEM[810];
assign MEM[2011] = MEM[306] + MEM[387];
assign MEM[2012] = MEM[309] + MEM[789];
assign MEM[2013] = MEM[311] + MEM[569];
assign MEM[2014] = MEM[314] + MEM[845];
assign MEM[2015] = MEM[316] + MEM[736];
assign MEM[2016] = MEM[316] + MEM[950];
assign MEM[2017] = MEM[317] + MEM[694];
assign MEM[2018] = MEM[318] + MEM[1280];
assign MEM[2019] = MEM[319] + MEM[1815];
assign MEM[2020] = MEM[322] + MEM[1110];
assign MEM[2021] = MEM[323] + MEM[480];
assign MEM[2022] = MEM[330] + MEM[918];
assign MEM[2023] = MEM[332] + MEM[1163];
assign MEM[2024] = MEM[336] + MEM[1026];
assign MEM[2025] = MEM[338] + MEM[1062];
assign MEM[2026] = MEM[339] + MEM[903];
assign MEM[2027] = MEM[341] + MEM[955];
assign MEM[2028] = MEM[342] + MEM[619];
assign MEM[2029] = MEM[350] + MEM[777];
assign MEM[2030] = MEM[354] + MEM[1100];
assign MEM[2031] = MEM[356] + MEM[359];
assign MEM[2032] = MEM[356] + MEM[683];
assign MEM[2033] = MEM[358] + MEM[747];
assign MEM[2034] = MEM[359] + MEM[1297];
assign MEM[2035] = MEM[362] + MEM[1027];
assign MEM[2036] = MEM[363] + MEM[398];
assign MEM[2037] = MEM[363] + MEM[1337];
assign MEM[2038] = MEM[364] + MEM[539];
assign MEM[2039] = MEM[370] + MEM[511];
assign MEM[2040] = MEM[370] + MEM[959];
assign MEM[2041] = MEM[371] + MEM[560];
assign MEM[2042] = MEM[371] + MEM[1008];
assign MEM[2043] = MEM[372] + MEM[526];
assign MEM[2044] = MEM[373] + MEM[602];
assign MEM[2045] = MEM[374] + MEM[761];
assign MEM[2046] = MEM[378] + MEM[940];
assign MEM[2047] = MEM[379] + MEM[1012];
assign MEM[2048] = MEM[380] + MEM[696];
assign MEM[2049] = MEM[380] + MEM[1135];
assign MEM[2050] = MEM[381] + MEM[805];
assign MEM[2051] = MEM[381] + MEM[812];
assign MEM[2052] = MEM[382] + MEM[415];
assign MEM[2053] = MEM[383] + MEM[421];
assign MEM[2054] = MEM[386] + MEM[1020];
assign MEM[2055] = MEM[388] + MEM[613];
assign MEM[2056] = MEM[389] + MEM[1331];
assign MEM[2057] = MEM[390] + MEM[915];
assign MEM[2058] = MEM[391] + MEM[834];
assign MEM[2059] = MEM[396] + MEM[466];
assign MEM[2060] = MEM[397] + MEM[1030];
assign MEM[2061] = MEM[399] + MEM[974];
assign MEM[2062] = MEM[403] + MEM[572];
assign MEM[2063] = MEM[406] + MEM[588];
assign MEM[2064] = MEM[410] + MEM[678];
assign MEM[2065] = MEM[412] + MEM[671];
assign MEM[2066] = MEM[414] + MEM[895];
assign MEM[2067] = MEM[416] + MEM[698];
assign MEM[2068] = MEM[417] + MEM[776];
assign MEM[2069] = MEM[421] + MEM[1194];
assign MEM[2070] = MEM[423] + MEM[498];
assign MEM[2071] = MEM[426] + MEM[715];
assign MEM[2072] = MEM[429] + MEM[1011];
assign MEM[2073] = MEM[430] + MEM[455];
assign MEM[2074] = MEM[431] + MEM[746];
assign MEM[2075] = MEM[435] + MEM[936];
assign MEM[2076] = MEM[436] + MEM[624];
assign MEM[2077] = MEM[438] + MEM[1167];
assign MEM[2078] = MEM[439] + MEM[1148];
assign MEM[2079] = MEM[439] + MEM[1263];
assign MEM[2080] = MEM[440] + MEM[698];
assign MEM[2081] = MEM[441] + MEM[690];
assign MEM[2082] = MEM[442] + MEM[900];
assign MEM[2083] = MEM[445] + MEM[1181];
assign MEM[2084] = MEM[448] + MEM[740];
assign MEM[2085] = MEM[449] + MEM[821];
assign MEM[2086] = MEM[451] + MEM[1350];
assign MEM[2087] = MEM[453] + MEM[1324];
assign MEM[2088] = MEM[454] + MEM[1156];
assign MEM[2089] = MEM[456] + MEM[705];
assign MEM[2090] = MEM[456] + MEM[1109];
assign MEM[2091] = MEM[457] + MEM[1088];
assign MEM[2092] = MEM[461] + MEM[1062];
assign MEM[2093] = MEM[462] + MEM[503];
assign MEM[2094] = MEM[464] + MEM[1632];
assign MEM[2095] = MEM[470] + MEM[819];
assign MEM[2096] = MEM[474] + MEM[947];
assign MEM[2097] = MEM[476] + MEM[652];
assign MEM[2098] = MEM[478] + MEM[1091];
assign MEM[2099] = MEM[482] + MEM[913];
assign MEM[2100] = MEM[483] + MEM[797];
assign MEM[2101] = MEM[485] + MEM[1133];
assign MEM[2102] = MEM[486] + MEM[825];
assign MEM[2103] = MEM[490] + MEM[689];
assign MEM[2104] = MEM[491] + MEM[804];
assign MEM[2105] = MEM[494] + MEM[979];
assign MEM[2106] = MEM[495] + MEM[599];
assign MEM[2107] = MEM[498] + MEM[1232];
assign MEM[2108] = MEM[513] + MEM[1391];
assign MEM[2109] = MEM[514] + MEM[837];
assign MEM[2110] = MEM[517] + MEM[800];
assign MEM[2111] = MEM[518] + MEM[1187];
assign MEM[2112] = MEM[519] + MEM[1518];
assign MEM[2113] = MEM[520] + MEM[958];
assign MEM[2114] = MEM[521] + MEM[1016];
assign MEM[2115] = MEM[524] + MEM[1676];
assign MEM[2116] = MEM[532] + MEM[1265];
assign MEM[2117] = MEM[540] + MEM[861];
assign MEM[2118] = MEM[541] + MEM[982];
assign MEM[2119] = MEM[544] + MEM[1532];
assign MEM[2120] = MEM[546] + MEM[565];
assign MEM[2121] = MEM[547] + MEM[573];
assign MEM[2122] = MEM[547] + MEM[660];
assign MEM[2123] = MEM[548] + MEM[761];
assign MEM[2124] = MEM[549] + MEM[1100];
assign MEM[2125] = MEM[552] + MEM[917];
assign MEM[2126] = MEM[556] + MEM[767];
assign MEM[2127] = MEM[558] + MEM[658];
assign MEM[2128] = MEM[559] + MEM[618];
assign MEM[2129] = MEM[561] + MEM[596];
assign MEM[2130] = MEM[564] + MEM[961];
assign MEM[2131] = MEM[566] + MEM[1184];
assign MEM[2132] = MEM[567] + MEM[593];
assign MEM[2133] = MEM[569] + MEM[625];
assign MEM[2134] = MEM[570] + MEM[1052];
assign MEM[2135] = MEM[571] + MEM[727];
assign MEM[2136] = MEM[573] + MEM[1196];
assign MEM[2137] = MEM[574] + MEM[863];
assign MEM[2138] = MEM[575] + MEM[870];
assign MEM[2139] = MEM[577] + MEM[796];
assign MEM[2140] = MEM[578] + MEM[632];
assign MEM[2141] = MEM[578] + MEM[1059];
assign MEM[2142] = MEM[581] + MEM[958];
assign MEM[2143] = MEM[584] + MEM[897];
assign MEM[2144] = MEM[587] + MEM[989];
assign MEM[2145] = MEM[589] + MEM[1146];
assign MEM[2146] = MEM[591] + MEM[672];
assign MEM[2147] = MEM[592] + MEM[749];
assign MEM[2148] = MEM[594] + MEM[704];
assign MEM[2149] = MEM[595] + MEM[633];
assign MEM[2150] = MEM[595] + MEM[1120];
assign MEM[2151] = MEM[596] + MEM[943];
assign MEM[2152] = MEM[597] + MEM[1050];
assign MEM[2153] = MEM[598] + MEM[989];
assign MEM[2154] = MEM[600] + MEM[925];
assign MEM[2155] = MEM[605] + MEM[752];
assign MEM[2156] = MEM[606] + MEM[1358];
assign MEM[2157] = MEM[607] + MEM[824];
assign MEM[2158] = MEM[609] + MEM[1004];
assign MEM[2159] = MEM[611] + MEM[695];
assign MEM[2160] = MEM[615] + MEM[994];
assign MEM[2161] = MEM[616] + MEM[1108];
assign MEM[2162] = MEM[620] + MEM[907];
assign MEM[2163] = MEM[621] + MEM[1544];
assign MEM[2164] = MEM[623] + MEM[780];
assign MEM[2165] = MEM[626] + MEM[914];
assign MEM[2166] = MEM[627] + MEM[1131];
assign MEM[2167] = MEM[628] + MEM[722];
assign MEM[2168] = MEM[629] + MEM[1189];
assign MEM[2169] = MEM[631] + MEM[1215];
assign MEM[2170] = MEM[632] + MEM[1253];
assign MEM[2171] = MEM[634] + MEM[901];
assign MEM[2172] = MEM[637] + MEM[1189];
assign MEM[2173] = MEM[638] + MEM[1705];
assign MEM[2174] = MEM[639] + MEM[1566];
assign MEM[2175] = MEM[645] + MEM[700];
assign MEM[2176] = MEM[646] + MEM[680];
assign MEM[2177] = MEM[648] + MEM[674];
assign MEM[2178] = MEM[649] + MEM[1069];
assign MEM[2179] = MEM[650] + MEM[1456];
assign MEM[2180] = MEM[652] + MEM[1210];
assign MEM[2181] = MEM[653] + MEM[787];
assign MEM[2182] = MEM[654] + MEM[656];
assign MEM[2183] = MEM[657] + MEM[1141];
assign MEM[2184] = MEM[659] + MEM[1146];
assign MEM[2185] = MEM[660] + MEM[1236];
assign MEM[2186] = MEM[661] + MEM[726];
assign MEM[2187] = MEM[662] + MEM[1545];
assign MEM[2188] = MEM[663] + MEM[708];
assign MEM[2189] = MEM[663] + MEM[1024];
assign MEM[2190] = MEM[664] + MEM[764];
assign MEM[2191] = MEM[665] + MEM[1326];
assign MEM[2192] = MEM[666] + MEM[876];
assign MEM[2193] = MEM[670] + MEM[1030];
assign MEM[2194] = MEM[672] + MEM[916];
assign MEM[2195] = MEM[673] + MEM[1043];
assign MEM[2196] = MEM[678] + MEM[868];
assign MEM[2197] = MEM[679] + MEM[855];
assign MEM[2198] = MEM[679] + MEM[1045];
assign MEM[2199] = MEM[680] + MEM[1066];
assign MEM[2200] = MEM[681] + MEM[722];
assign MEM[2201] = MEM[683] + MEM[906];
assign MEM[2202] = MEM[684] + MEM[969];
assign MEM[2203] = MEM[685] + MEM[1079];
assign MEM[2204] = MEM[688] + MEM[1082];
assign MEM[2205] = MEM[693] + MEM[769];
assign MEM[2206] = MEM[693] + MEM[1118];
assign MEM[2207] = MEM[694] + MEM[789];
assign MEM[2208] = MEM[697] + MEM[1303];
assign MEM[2209] = MEM[699] + MEM[1044];
assign MEM[2210] = MEM[702] + MEM[1264];
assign MEM[2211] = MEM[703] + MEM[1344];
assign MEM[2212] = MEM[706] + MEM[959];
assign MEM[2213] = MEM[710] + MEM[838];
assign MEM[2214] = MEM[711] + MEM[784];
assign MEM[2215] = MEM[711] + MEM[887];
assign MEM[2216] = MEM[713] + MEM[1278];
assign MEM[2217] = MEM[714] + MEM[740];
assign MEM[2218] = MEM[716] + MEM[743];
assign MEM[2219] = MEM[719] + MEM[1147];
assign MEM[2220] = MEM[720] + MEM[881];
assign MEM[2221] = MEM[723] + MEM[1027];
assign MEM[2222] = MEM[734] + MEM[782];
assign MEM[2223] = MEM[735] + MEM[1101];
assign MEM[2224] = MEM[736] + MEM[954];
assign MEM[2225] = MEM[737] + MEM[1182];
assign MEM[2226] = MEM[738] + MEM[1207];
assign MEM[2227] = MEM[741] + MEM[1072];
assign MEM[2228] = MEM[742] + MEM[1143];
assign MEM[2229] = MEM[744] + MEM[1323];
assign MEM[2230] = MEM[745] + MEM[1034];
assign MEM[2231] = MEM[747] + MEM[1085];
assign MEM[2232] = MEM[748] + MEM[1311];
assign MEM[2233] = MEM[752] + MEM[993];
assign MEM[2234] = MEM[755] + MEM[960];
assign MEM[2235] = MEM[758] + MEM[1172];
assign MEM[2236] = MEM[759] + MEM[1199];
assign MEM[2237] = MEM[760] + MEM[1157];
assign MEM[2238] = MEM[763] + MEM[848];
assign MEM[2239] = MEM[764] + MEM[1067];
assign MEM[2240] = MEM[765] + MEM[1089];
assign MEM[2241] = MEM[768] + MEM[1295];
assign MEM[2242] = MEM[771] + MEM[1152];
assign MEM[2243] = MEM[772] + MEM[1208];
assign MEM[2244] = MEM[773] + MEM[923];
assign MEM[2245] = MEM[774] + MEM[2062];
assign MEM[2246] = MEM[775] + MEM[902];
assign MEM[2247] = MEM[778] + MEM[1596];
assign MEM[2248] = MEM[779] + MEM[1283];
assign MEM[2249] = MEM[780] + MEM[1200];
assign MEM[2250] = MEM[783] + MEM[873];
assign MEM[2251] = MEM[786] + MEM[1333];
assign MEM[2252] = MEM[787] + MEM[877];
assign MEM[2253] = MEM[788] + MEM[1143];
assign MEM[2254] = MEM[790] + MEM[886];
assign MEM[2255] = MEM[793] + MEM[845];
assign MEM[2256] = MEM[794] + MEM[840];
assign MEM[2257] = MEM[795] + MEM[1080];
assign MEM[2258] = MEM[796] + MEM[1072];
assign MEM[2259] = MEM[798] + MEM[1217];
assign MEM[2260] = MEM[799] + MEM[1464];
assign MEM[2261] = MEM[800] + MEM[1418];
assign MEM[2262] = MEM[802] + MEM[936];
assign MEM[2263] = MEM[803] + MEM[1219];
assign MEM[2264] = MEM[806] + MEM[1243];
assign MEM[2265] = MEM[808] + MEM[1082];
assign MEM[2266] = MEM[808] + MEM[1573];
assign MEM[2267] = MEM[809] + MEM[959];
assign MEM[2268] = MEM[812] + MEM[1299];
assign MEM[2269] = MEM[813] + MEM[1041];
assign MEM[2270] = MEM[816] + MEM[1125];
assign MEM[2271] = MEM[817] + MEM[909];
assign MEM[2272] = MEM[818] + MEM[1804];
assign MEM[2273] = MEM[819] + MEM[1081];
assign MEM[2274] = MEM[820] + MEM[831];
assign MEM[2275] = MEM[823] + MEM[1040];
assign MEM[2276] = MEM[827] + MEM[885];
assign MEM[2277] = MEM[828] + MEM[1459];
assign MEM[2278] = MEM[829] + MEM[1017];
assign MEM[2279] = MEM[830] + MEM[1089];
assign MEM[2280] = MEM[831] + MEM[839];
assign MEM[2281] = MEM[832] + MEM[1375];
assign MEM[2282] = MEM[834] + MEM[974];
assign MEM[2283] = MEM[834] + MEM[1405];
assign MEM[2284] = MEM[835] + MEM[983];
assign MEM[2285] = MEM[836] + MEM[920];
assign MEM[2286] = MEM[838] + MEM[1949];
assign MEM[2287] = MEM[839] + MEM[1123];
assign MEM[2288] = MEM[840] + MEM[1004];
assign MEM[2289] = MEM[841] + MEM[968];
assign MEM[2290] = MEM[843] + MEM[942];
assign MEM[2291] = MEM[844] + MEM[1036];
assign MEM[2292] = MEM[845] + MEM[1477];
assign MEM[2293] = MEM[846] + MEM[1302];
assign MEM[2294] = MEM[847] + MEM[952];
assign MEM[2295] = MEM[847] + MEM[981];
assign MEM[2296] = MEM[850] + MEM[866];
assign MEM[2297] = MEM[851] + MEM[996];
assign MEM[2298] = MEM[853] + MEM[924];
assign MEM[2299] = MEM[853] + MEM[1292];
assign MEM[2300] = MEM[854] + MEM[1436];
assign MEM[2301] = MEM[856] + MEM[1106];
assign MEM[2302] = MEM[857] + MEM[1118];
assign MEM[2303] = MEM[858] + MEM[1058];
assign MEM[2304] = MEM[859] + MEM[934];
assign MEM[2305] = MEM[860] + MEM[1208];
assign MEM[2306] = MEM[864] + MEM[1114];
assign MEM[2307] = MEM[867] + MEM[1221];
assign MEM[2308] = MEM[869] + MEM[1169];
assign MEM[2309] = MEM[870] + MEM[1313];
assign MEM[2310] = MEM[871] + MEM[935];
assign MEM[2311] = MEM[873] + MEM[1110];
assign MEM[2312] = MEM[874] + MEM[1003];
assign MEM[2313] = MEM[875] + MEM[1183];
assign MEM[2314] = MEM[877] + MEM[1344];
assign MEM[2315] = MEM[879] + MEM[1542];
assign MEM[2316] = MEM[881] + MEM[1028];
assign MEM[2317] = MEM[883] + MEM[1700];
assign MEM[2318] = MEM[885] + MEM[1266];
assign MEM[2319] = MEM[888] + MEM[1075];
assign MEM[2320] = MEM[891] + MEM[1198];
assign MEM[2321] = MEM[892] + MEM[1332];
assign MEM[2322] = MEM[893] + MEM[1095];
assign MEM[2323] = MEM[894] + MEM[1404];
assign MEM[2324] = MEM[896] + MEM[953];
assign MEM[2325] = MEM[896] + MEM[1222];
assign MEM[2326] = MEM[897] + MEM[1137];
assign MEM[2327] = MEM[898] + MEM[985];
assign MEM[2328] = MEM[898] + MEM[1179];
assign MEM[2329] = MEM[899] + MEM[1363];
assign MEM[2330] = MEM[900] + MEM[1342];
assign MEM[2331] = MEM[902] + MEM[1074];
assign MEM[2332] = MEM[903] + MEM[1188];
assign MEM[2333] = MEM[906] + MEM[1587];
assign MEM[2334] = MEM[908] + MEM[1187];
assign MEM[2335] = MEM[910] + MEM[990];
assign MEM[2336] = MEM[912] + MEM[1610];
assign MEM[2337] = MEM[914] + MEM[1028];
assign MEM[2338] = MEM[916] + MEM[1251];
assign MEM[2339] = MEM[917] + MEM[1280];
assign MEM[2340] = MEM[918] + MEM[1068];
assign MEM[2341] = MEM[924] + MEM[1600];
assign MEM[2342] = MEM[925] + MEM[1017];
assign MEM[2343] = MEM[928] + MEM[1056];
assign MEM[2344] = MEM[928] + MEM[1538];
assign MEM[2345] = MEM[931] + MEM[1695];
assign MEM[2346] = MEM[934] + MEM[1261];
assign MEM[2347] = MEM[935] + MEM[1467];
assign MEM[2348] = MEM[940] + MEM[1215];
assign MEM[2349] = MEM[941] + MEM[1088];
assign MEM[2350] = MEM[942] + MEM[1389];
assign MEM[2351] = MEM[944] + MEM[1119];
assign MEM[2352] = MEM[945] + MEM[1052];
assign MEM[2353] = MEM[947] + MEM[1279];
assign MEM[2354] = MEM[948] + MEM[1334];
assign MEM[2355] = MEM[950] + MEM[1180];
assign MEM[2356] = MEM[952] + MEM[1240];
assign MEM[2357] = MEM[953] + MEM[1175];
assign MEM[2358] = MEM[954] + MEM[1252];
assign MEM[2359] = MEM[955] + MEM[1657];
assign MEM[2360] = MEM[956] + MEM[1296];
assign MEM[2361] = MEM[957] + MEM[1027];
assign MEM[2362] = MEM[962] + MEM[1209];
assign MEM[2363] = MEM[964] + MEM[1018];
assign MEM[2364] = MEM[965] + MEM[1178];
assign MEM[2365] = MEM[966] + MEM[976];
assign MEM[2366] = MEM[967] + MEM[1268];
assign MEM[2367] = MEM[973] + MEM[1055];
assign MEM[2368] = MEM[974] + MEM[1201];
assign MEM[2369] = MEM[975] + MEM[1127];
assign MEM[2370] = MEM[977] + MEM[1134];
assign MEM[2371] = MEM[978] + MEM[1007];
assign MEM[2372] = MEM[980] + MEM[1049];
assign MEM[2373] = MEM[982] + MEM[1120];
assign MEM[2374] = MEM[984] + MEM[1353];
assign MEM[2375] = MEM[987] + MEM[1369];
assign MEM[2376] = MEM[988] + MEM[1216];
assign MEM[2377] = MEM[989] + MEM[1200];
assign MEM[2378] = MEM[992] + MEM[1126];
assign MEM[2379] = MEM[995] + MEM[1158];
assign MEM[2380] = MEM[997] + MEM[1000];
assign MEM[2381] = MEM[999] + MEM[1019];
assign MEM[2382] = MEM[1001] + MEM[1129];
assign MEM[2383] = MEM[1004] + MEM[1317];
assign MEM[2384] = MEM[1005] + MEM[1332];
assign MEM[2385] = MEM[1012] + MEM[1103];
assign MEM[2386] = MEM[1012] + MEM[1799];
assign MEM[2387] = MEM[1013] + MEM[1099];
assign MEM[2388] = MEM[1015] + MEM[1321];
assign MEM[2389] = MEM[1017] + MEM[1284];
assign MEM[2390] = MEM[1018] + MEM[1236];
assign MEM[2391] = MEM[1020] + MEM[1047];
assign MEM[2392] = MEM[1020] + MEM[1489];
assign MEM[2393] = MEM[1021] + MEM[1340];
assign MEM[2394] = MEM[1022] + MEM[1204];
assign MEM[2395] = MEM[1023] + MEM[1756];
assign MEM[2396] = MEM[1028] + MEM[1584];
assign MEM[2397] = MEM[1031] + MEM[1310];
assign MEM[2398] = MEM[1032] + MEM[1051];
assign MEM[2399] = MEM[1035] + MEM[1102];
assign MEM[2400] = MEM[1038] + MEM[1119];
assign MEM[2401] = MEM[1039] + MEM[1371];
assign MEM[2402] = MEM[1046] + MEM[1079];
assign MEM[2403] = MEM[1057] + MEM[1621];
assign MEM[2404] = MEM[1058] + MEM[1097];
assign MEM[2405] = MEM[1058] + MEM[1309];
assign MEM[2406] = MEM[1060] + MEM[1177];
assign MEM[2407] = MEM[1061] + MEM[1347];
assign MEM[2408] = MEM[1062] + MEM[1186];
assign MEM[2409] = MEM[1063] + MEM[1095];
assign MEM[2410] = MEM[1065] + MEM[1202];
assign MEM[2411] = MEM[1066] + MEM[1310];
assign MEM[2412] = MEM[1069] + MEM[1109];
assign MEM[2413] = MEM[1069] + MEM[1195];
assign MEM[2414] = MEM[1070] + MEM[1223];
assign MEM[2415] = MEM[1073] + MEM[1279];
assign MEM[2416] = MEM[1074] + MEM[1411];
assign MEM[2417] = MEM[1076] + MEM[1514];
assign MEM[2418] = MEM[1077] + MEM[1362];
assign MEM[2419] = MEM[1080] + MEM[1491];
assign MEM[2420] = MEM[1083] + MEM[1195];
assign MEM[2421] = MEM[1083] + MEM[1673];
assign MEM[2422] = MEM[1084] + MEM[1273];
assign MEM[2423] = MEM[1085] + MEM[1127];
assign MEM[2424] = MEM[1086] + MEM[1278];
assign MEM[2425] = MEM[1087] + MEM[1325];
assign MEM[2426] = MEM[1090] + MEM[2015];
assign MEM[2427] = MEM[1091] + MEM[1205];
assign MEM[2428] = MEM[1092] + MEM[1468];
assign MEM[2429] = MEM[1093] + MEM[1356];
assign MEM[2430] = MEM[1094] + MEM[1458];
assign MEM[2431] = MEM[1096] + MEM[1382];
assign MEM[2432] = MEM[1098] + MEM[1305];
assign MEM[2433] = MEM[1099] + MEM[1524];
assign MEM[2434] = MEM[1102] + MEM[1103];
assign MEM[2435] = MEM[1104] + MEM[1214];
assign MEM[2436] = MEM[1105] + MEM[1287];
assign MEM[2437] = MEM[1107] + MEM[1618];
assign MEM[2438] = MEM[1111] + MEM[1366];
assign MEM[2439] = MEM[1112] + MEM[1154];
assign MEM[2440] = MEM[1113] + MEM[1486];
assign MEM[2441] = MEM[1115] + MEM[1291];
assign MEM[2442] = MEM[1116] + MEM[1306];
assign MEM[2443] = MEM[1117] + MEM[1177];
assign MEM[2444] = MEM[1121] + MEM[1288];
assign MEM[2445] = MEM[1124] + MEM[1173];
assign MEM[2446] = MEM[1126] + MEM[1163];
assign MEM[2447] = MEM[1129] + MEM[1211];
assign MEM[2448] = MEM[1132] + MEM[1959];
assign MEM[2449] = MEM[1133] + MEM[1269];
assign MEM[2450] = MEM[1135] + MEM[1761];
assign MEM[2451] = MEM[1136] + MEM[1273];
assign MEM[2452] = MEM[1137] + MEM[1388];
assign MEM[2453] = MEM[1138] + MEM[1655];
assign MEM[2454] = MEM[1139] + MEM[1266];
assign MEM[2455] = MEM[1140] + MEM[2121];
assign MEM[2456] = MEM[1141] + MEM[1424];
assign MEM[2457] = MEM[1142] + MEM[1284];
assign MEM[2458] = MEM[1144] + MEM[1222];
assign MEM[2459] = MEM[1145] + MEM[1678];
assign MEM[2460] = MEM[1147] + MEM[1196];
assign MEM[2461] = MEM[1148] + MEM[1167];
assign MEM[2462] = MEM[1149] + MEM[1312];
assign MEM[2463] = MEM[1150] + MEM[1560];
assign MEM[2464] = MEM[1153] + MEM[1134];
assign MEM[2465] = MEM[1154] + MEM[1218];
assign MEM[2466] = MEM[1157] + MEM[1250];
assign MEM[2467] = MEM[1158] + MEM[1461];
assign MEM[2468] = MEM[1159] + MEM[1419];
assign MEM[2469] = MEM[1160] + MEM[1585];
assign MEM[2470] = MEM[1161] + MEM[1329];
assign MEM[2471] = MEM[1162] + MEM[1245];
assign MEM[2472] = MEM[1162] + MEM[1248];
assign MEM[2473] = MEM[1164] + MEM[1443];
assign MEM[2474] = MEM[1165] + MEM[1270];
assign MEM[2475] = MEM[1165] + MEM[1286];
assign MEM[2476] = MEM[1166] + MEM[2398];
assign MEM[2477] = MEM[1168] + MEM[1743];
assign MEM[2478] = MEM[1169] + MEM[1408];
assign MEM[2479] = MEM[1170] + MEM[1292];
assign MEM[2480] = MEM[1171] + MEM[1691];
assign MEM[2481] = MEM[1172] + MEM[1225];
assign MEM[2482] = MEM[1174] + MEM[1696];
assign MEM[2483] = MEM[1175] + MEM[1370];
assign MEM[2484] = MEM[1176] + MEM[1475];
assign MEM[2485] = MEM[1179] + MEM[1694];
assign MEM[2486] = MEM[1181] + MEM[1228];
assign MEM[2487] = MEM[1184] + MEM[1341];
assign MEM[2488] = MEM[1185] + MEM[1247];
assign MEM[2489] = MEM[1190] + MEM[1470];
assign MEM[2490] = MEM[1191] + MEM[1256];
assign MEM[2491] = MEM[1192] + MEM[1293];
assign MEM[2492] = MEM[1197] + MEM[1326];
assign MEM[2493] = MEM[1197] + MEM[1397];
assign MEM[2494] = MEM[1202] + MEM[1226];
assign MEM[2495] = MEM[1204] + MEM[1738];
assign MEM[2496] = MEM[1205] + MEM[1212];
assign MEM[2497] = MEM[1206] + MEM[1277];
assign MEM[2498] = MEM[1206] + MEM[1472];
assign MEM[2499] = MEM[1207] + MEM[1314];
assign MEM[2500] = MEM[1209] + MEM[1380];
assign MEM[2501] = MEM[1210] + MEM[1481];
assign MEM[2502] = MEM[1211] + MEM[1328];
assign MEM[2503] = MEM[1213] + MEM[1364];
assign MEM[2504] = MEM[1214] + MEM[1772];
assign MEM[2505] = MEM[1216] + MEM[1499];
assign MEM[2506] = MEM[1217] + MEM[1437];
assign MEM[2507] = MEM[1218] + MEM[1619];
assign MEM[2508] = MEM[1219] + MEM[1564];
assign MEM[2509] = MEM[1220] + MEM[1563];
assign MEM[2510] = MEM[1223] + MEM[1415];
assign MEM[2511] = MEM[1224] + MEM[2133];
assign MEM[2512] = MEM[1225] + MEM[1241];
assign MEM[2513] = MEM[1227] + MEM[1246];
assign MEM[2514] = MEM[1229] + MEM[1304];
assign MEM[2515] = MEM[1231] + MEM[1692];
assign MEM[2516] = MEM[1232] + MEM[1728];
assign MEM[2517] = MEM[1234] + MEM[1614];
assign MEM[2518] = MEM[1234] + MEM[2445];
assign MEM[2519] = MEM[1235] + MEM[1455];
assign MEM[2520] = MEM[1238] + MEM[1327];
assign MEM[2521] = MEM[1238] + MEM[1599];
assign MEM[2522] = MEM[1239] + MEM[1633];
assign MEM[2523] = MEM[1240] + MEM[1435];
assign MEM[2524] = MEM[1242] + MEM[1346];
assign MEM[2525] = MEM[1243] + MEM[1495];
assign MEM[2526] = MEM[1244] + MEM[1307];
assign MEM[2527] = MEM[1244] + MEM[1333];
assign MEM[2528] = MEM[1246] + MEM[1505];
assign MEM[2529] = MEM[1247] + MEM[1249];
assign MEM[2530] = MEM[1248] + MEM[1315];
assign MEM[2531] = MEM[1250] + MEM[1429];
assign MEM[2532] = MEM[1252] + MEM[1604];
assign MEM[2533] = MEM[1253] + MEM[1745];
assign MEM[2534] = MEM[1254] + MEM[849];
assign MEM[2535] = MEM[1257] + MEM[1271];
assign MEM[2536] = MEM[1257] + MEM[1767];
assign MEM[2537] = MEM[1258] + MEM[1448];
assign MEM[2538] = MEM[1258] + MEM[1675];
assign MEM[2539] = MEM[1260] + MEM[1272];
assign MEM[2540] = MEM[1261] + MEM[1697];
assign MEM[2541] = MEM[1262] + MEM[1629];
assign MEM[2542] = MEM[1262] + MEM[1941];
assign MEM[2543] = MEM[1264] + MEM[1506];
assign MEM[2544] = MEM[1267] + MEM[1311];
assign MEM[2545] = MEM[1268] + MEM[2376];
assign MEM[2546] = MEM[1271] + MEM[1658];
assign MEM[2547] = MEM[1274] + MEM[1541];
assign MEM[2548] = MEM[1276] + MEM[1335];
assign MEM[2549] = MEM[1276] + MEM[1452];
assign MEM[2550] = MEM[1281] + MEM[1308];
assign MEM[2551] = MEM[1281] + MEM[1942];
assign MEM[2552] = MEM[1282] + MEM[1662];
assign MEM[2553] = MEM[1282] + MEM[1748];
assign MEM[2554] = MEM[1285] + MEM[1329];
assign MEM[2555] = MEM[1285] + MEM[2220];
assign MEM[2556] = MEM[1287] + MEM[1352];
assign MEM[2557] = MEM[1289] + MEM[2423];
assign MEM[2558] = MEM[1290] + MEM[1354];
assign MEM[2559] = MEM[1293] + MEM[1392];
assign MEM[2560] = MEM[1294] + MEM[1357];
assign MEM[2561] = MEM[1294] + MEM[1620];
assign MEM[2562] = MEM[1295] + MEM[2287];
assign MEM[2563] = MEM[1299] + MEM[1351];
assign MEM[2564] = MEM[1301] + MEM[1719];
assign MEM[2565] = MEM[1302] + MEM[1634];
assign MEM[2566] = MEM[1303] + MEM[2296];
assign MEM[2567] = MEM[1304] + MEM[1438];
assign MEM[2568] = MEM[1305] + MEM[1715];
assign MEM[2569] = MEM[1306] + MEM[1623];
assign MEM[2570] = MEM[1307] + MEM[1591];
assign MEM[2571] = MEM[1309] + MEM[2182];
assign MEM[2572] = MEM[1312] + MEM[1725];
assign MEM[2573] = MEM[1313] + MEM[1654];
assign MEM[2574] = MEM[1314] + MEM[1746];
assign MEM[2575] = MEM[1315] + MEM[1422];
assign MEM[2576] = MEM[1318] + MEM[1361];
assign MEM[2577] = MEM[1319] + MEM[1423];
assign MEM[2578] = MEM[1319] + MEM[1636];
assign MEM[2579] = MEM[1320] + MEM[1450];
assign MEM[2580] = MEM[1320] + MEM[1641];
assign MEM[2581] = MEM[1321] + MEM[1553];
assign MEM[2582] = MEM[1322] + MEM[1447];
assign MEM[2583] = MEM[1322] + MEM[1469];
assign MEM[2584] = MEM[1323] + MEM[1707];
assign MEM[2585] = MEM[1325] + MEM[1583];
assign MEM[2586] = MEM[1327] + MEM[2071];
assign MEM[2587] = MEM[1328] + MEM[1708];
assign MEM[2588] = MEM[1330] + MEM[1433];
assign MEM[2589] = MEM[1330] + MEM[1921];
assign MEM[2590] = MEM[1334] + MEM[2409];
assign MEM[2591] = MEM[1335] + MEM[1607];
assign MEM[2592] = MEM[1336] + MEM[1478];
assign MEM[2593] = MEM[1336] + MEM[1565];
assign MEM[2594] = MEM[1338] + MEM[1364];
assign MEM[2595] = MEM[1338] + MEM[2197];
assign MEM[2596] = MEM[1339] + MEM[1390];
assign MEM[2597] = MEM[1339] + MEM[1773];
assign MEM[2598] = MEM[1340] + MEM[1740];
assign MEM[2599] = MEM[1343] + MEM[1465];
assign MEM[2600] = MEM[1345] + MEM[1454];
assign MEM[2601] = MEM[1345] + MEM[1581];
assign MEM[2602] = MEM[1347] + MEM[1387];
assign MEM[2603] = MEM[1348] + MEM[1690];
assign MEM[2604] = MEM[1349] + MEM[1373];
assign MEM[2605] = MEM[1351] + MEM[1612];
assign MEM[2606] = MEM[1352] + MEM[1552];
assign MEM[2607] = MEM[1353] + MEM[1403];
assign MEM[2608] = MEM[1354] + MEM[1859];
assign MEM[2609] = MEM[1355] + MEM[1360];
assign MEM[2610] = MEM[1355] + MEM[1782];
assign MEM[2611] = MEM[1356] + MEM[1551];
assign MEM[2612] = MEM[1357] + MEM[1471];
assign MEM[2613] = MEM[1359] + MEM[1543];
assign MEM[2614] = MEM[1360] + MEM[2167];
assign MEM[2615] = MEM[1362] + MEM[1681];
assign MEM[2616] = MEM[1363] + MEM[1558];
assign MEM[2617] = MEM[1365] + MEM[1523];
assign MEM[2618] = MEM[1368] + MEM[1485];
assign MEM[2619] = MEM[1369] + MEM[1384];
assign MEM[2620] = MEM[1371] + MEM[2134];
assign MEM[2621] = MEM[1372] + MEM[1513];
assign MEM[2622] = MEM[1372] + MEM[1660];
assign MEM[2623] = MEM[1374] + MEM[1421];
assign MEM[2624] = MEM[1374] + MEM[1439];
assign MEM[2625] = MEM[1375] + MEM[1378];
assign MEM[2626] = MEM[1377] + MEM[1530];
assign MEM[2627] = MEM[1379] + MEM[1734];
assign MEM[2628] = MEM[1381] + MEM[2107];
assign MEM[2629] = MEM[1385] + MEM[1789];
assign MEM[2630] = MEM[1393] + MEM[1645];
assign MEM[2631] = MEM[1394] + MEM[1383];
assign MEM[2632] = MEM[1395] + MEM[1651];
assign MEM[2633] = MEM[1398] + MEM[1605];
assign MEM[2634] = MEM[1399] + MEM[1504];
assign MEM[2635] = MEM[1400] + MEM[1401];
assign MEM[2636] = MEM[1410] + MEM[1511];
assign MEM[2637] = MEM[1413] + MEM[1597];
assign MEM[2638] = MEM[1414] + MEM[2068];
assign MEM[2639] = MEM[1416] + MEM[1689];
assign MEM[2640] = MEM[1425] + MEM[1578];
assign MEM[2641] = MEM[1426] + MEM[2122];
assign MEM[2642] = MEM[1427] + MEM[1908];
assign MEM[2643] = MEM[1428] + MEM[1582];
assign MEM[2644] = MEM[1430] + MEM[1457];
assign MEM[2645] = MEM[1434] + MEM[2089];
assign MEM[2646] = MEM[1440] + MEM[1763];
assign MEM[2647] = MEM[1446] + MEM[1814];
assign MEM[2648] = MEM[1449] + MEM[1751];
assign MEM[2649] = MEM[1451] + MEM[1115];
assign MEM[2650] = MEM[1453] + MEM[1753];
assign MEM[2651] = MEM[1460] + MEM[1586];
assign MEM[2652] = MEM[1473] + MEM[1482];
assign MEM[2653] = MEM[1474] + MEM[1682];
assign MEM[2654] = MEM[1483] + MEM[1724];
assign MEM[2655] = MEM[1484] + MEM[1527];
assign MEM[2656] = MEM[1487] + MEM[1648];
assign MEM[2657] = MEM[1488] + MEM[1556];
assign MEM[2658] = MEM[1492] + MEM[1752];
assign MEM[2659] = MEM[1494] + MEM[1788];
assign MEM[2660] = MEM[1496] + MEM[1512];
assign MEM[2661] = MEM[1497] + MEM[1649];
assign MEM[2662] = MEM[1498] + MEM[1887];
assign MEM[2663] = MEM[1500] + MEM[1754];
assign MEM[2664] = MEM[1502] + MEM[1576];
assign MEM[2665] = MEM[1507] + MEM[1741];
assign MEM[2666] = MEM[1508] + MEM[1744];
assign MEM[2667] = MEM[1509] + MEM[1517];
assign MEM[2668] = MEM[1516] + MEM[1861];
assign MEM[2669] = MEM[1519] + MEM[1812];
assign MEM[2670] = MEM[1520] + MEM[1562];
assign MEM[2671] = MEM[1521] + MEM[1727];
assign MEM[2672] = MEM[1522] + MEM[1550];
assign MEM[2673] = MEM[1525] + MEM[1793];
assign MEM[2674] = MEM[1526] + MEM[1800];
assign MEM[2675] = MEM[1528] + MEM[1731];
assign MEM[2676] = MEM[1529] + MEM[1592];
assign MEM[2677] = MEM[1531] + MEM[1630];
assign MEM[2678] = MEM[1537] + MEM[2085];
assign MEM[2679] = MEM[1548] + MEM[1669];
assign MEM[2680] = MEM[1554] + MEM[1653];
assign MEM[2681] = MEM[1555] + MEM[1547];
assign MEM[2682] = MEM[1561] + MEM[1693];
assign MEM[2683] = MEM[1569] + MEM[2084];
assign MEM[2684] = MEM[1570] + MEM[2506];
assign MEM[2685] = MEM[1571] + MEM[1980];
assign MEM[2686] = MEM[1572] + MEM[1764];
assign MEM[2687] = MEM[1574] + MEM[1755];
assign MEM[2688] = MEM[1575] + MEM[1983];
assign MEM[2689] = MEM[1579] + MEM[1713];
assign MEM[2690] = MEM[1580] + MEM[1801];
assign MEM[2691] = MEM[1588] + MEM[2229];
assign MEM[2692] = MEM[1589] + MEM[1602];
assign MEM[2693] = MEM[1590] + MEM[1515];
assign MEM[2694] = MEM[1594] + MEM[1795];
assign MEM[2695] = MEM[1601] + MEM[1650];
assign MEM[2696] = MEM[1603] + MEM[1779];
assign MEM[2697] = MEM[1608] + MEM[2396];
assign MEM[2698] = MEM[1611] + MEM[1656];
assign MEM[2699] = MEM[1616] + MEM[1642];
assign MEM[2700] = MEM[1624] + MEM[1652];
assign MEM[2701] = MEM[1631] + MEM[2034];
assign MEM[2702] = MEM[1638] + MEM[1199];
assign MEM[2703] = MEM[1643] + MEM[1994];
assign MEM[2704] = MEM[1646] + MEM[1762];
assign MEM[2705] = MEM[1647] + MEM[1701];
assign MEM[2706] = MEM[1659] + MEM[1784];
assign MEM[2707] = MEM[1661] + MEM[1714];
assign MEM[2708] = MEM[1668] + MEM[1683];
assign MEM[2709] = MEM[1679] + MEM[2494];
assign MEM[2710] = MEM[1685] + MEM[1759];
assign MEM[2711] = MEM[1687] + MEM[1839];
assign MEM[2712] = MEM[1688] + MEM[1771];
assign MEM[2713] = MEM[1698] + MEM[1720];
assign MEM[2714] = MEM[1703] + MEM[2268];
assign MEM[2715] = MEM[1709] + MEM[2011];
assign MEM[2716] = MEM[1712] + MEM[1717];
assign MEM[2717] = MEM[1716] + MEM[1913];
assign MEM[2718] = MEM[1721] + MEM[1723];
assign MEM[2719] = MEM[1722] + MEM[1910];
assign MEM[2720] = MEM[1730] + MEM[2004];
assign MEM[2721] = MEM[1742] + MEM[1819];
assign MEM[2722] = MEM[1749] + MEM[2322];
assign MEM[2723] = MEM[1750] + MEM[1857];
assign MEM[2724] = MEM[1758] + MEM[1955];
assign MEM[2725] = MEM[1783] + MEM[2527];
assign MEM[2726] = MEM[1794] + MEM[2169];
assign MEM[2727] = MEM[1796] + MEM[2211];
assign MEM[2728] = MEM[1805] + MEM[1832];
assign MEM[2729] = MEM[1808] + MEM[1823];
assign MEM[2730] = MEM[1810] + MEM[1830];
assign MEM[2731] = MEM[1811] + MEM[1536];
assign MEM[2732] = MEM[1833] + MEM[2316];
assign MEM[2733] = MEM[1843] + MEM[2530];
assign MEM[2734] = MEM[1844] + MEM[2400];
assign MEM[2735] = MEM[1848] + MEM[1792];
assign MEM[2736] = MEM[1849] + MEM[2261];
assign MEM[2737] = MEM[1850] + MEM[2611];
assign MEM[2738] = MEM[1851] + MEM[2501];
assign MEM[2739] = MEM[1852] + MEM[2399];
assign MEM[2740] = MEM[1853] + MEM[2353];
assign MEM[2741] = MEM[1863] + MEM[2609];
assign MEM[2742] = MEM[1864] + MEM[1786];
assign MEM[2743] = MEM[1869] + MEM[1670];
assign MEM[2744] = MEM[1870] + MEM[1798];
assign MEM[2745] = MEM[1872] + MEM[1677];
assign MEM[2746] = MEM[1876] + MEM[2054];
assign MEM[2747] = MEM[1891] + MEM[2480];
assign MEM[2748] = MEM[1909] + MEM[2513];
assign MEM[2749] = MEM[1911] + MEM[2368];
assign MEM[2750] = MEM[1914] + MEM[2622];
assign MEM[2751] = MEM[1916] + MEM[2161];
assign MEM[2752] = MEM[1917] + MEM[1640];
assign MEM[2753] = MEM[1918] + MEM[1615];
assign MEM[2754] = MEM[1923] + MEM[2114];
assign MEM[2755] = MEM[1924] + MEM[2559];
assign MEM[2756] = MEM[1926] + MEM[2643];
assign MEM[2757] = MEM[1930] + MEM[2629];
assign MEM[2758] = MEM[1931] + MEM[2140];
assign MEM[2759] = MEM[1934] + MEM[1726];
assign MEM[2760] = MEM[1937] + MEM[2408];
assign MEM[2761] = MEM[1940] + MEM[2615];
assign MEM[2762] = MEM[1945] + MEM[2627];
assign MEM[2763] = MEM[1954] + MEM[2305];
assign MEM[2764] = MEM[1960] + MEM[2516];
assign MEM[2765] = MEM[1963] + MEM[2326];
assign MEM[2766] = MEM[1965] + MEM[2246];
assign MEM[2767] = MEM[1972] + MEM[2435];
assign MEM[2768] = MEM[1974] + MEM[2630];
assign MEM[2769] = MEM[1979] + MEM[2152];
assign MEM[2770] = MEM[1981] + MEM[2547];
assign MEM[2771] = MEM[1982] + MEM[2694];
assign MEM[2772] = MEM[1984] + MEM[2531];
assign MEM[2773] = MEM[1989] + MEM[1775];
assign MEM[2774] = MEM[1997] + MEM[2477];
assign MEM[2775] = MEM[2002] + MEM[2544];
assign MEM[2776] = MEM[2005] + MEM[2673];
assign MEM[2777] = MEM[2006] + MEM[2648];
assign MEM[2778] = MEM[2013] + MEM[2165];
assign MEM[2779] = MEM[2025] + MEM[2695];
assign MEM[2780] = MEM[2026] + MEM[2660];
assign MEM[2781] = MEM[2029] + MEM[2249];
assign MEM[2782] = MEM[2036] + MEM[2079];
assign MEM[2783] = MEM[2039] + MEM[2116];
assign MEM[2784] = MEM[2040] + MEM[2657];
assign MEM[2785] = MEM[2041] + MEM[2427];
assign MEM[2786] = MEM[2042] + MEM[1666];
assign MEM[2787] = MEM[2043] + MEM[2446];
assign MEM[2788] = MEM[2044] + MEM[2686];
assign MEM[2789] = MEM[2049] + MEM[2505];
assign MEM[2790] = MEM[2050] + MEM[2700];
assign MEM[2791] = MEM[2053] + MEM[2073];
assign MEM[2792] = MEM[2055] + MEM[2251];
assign MEM[2793] = MEM[2057] + MEM[2416];
assign MEM[2794] = MEM[2083] + MEM[2689];
assign MEM[2795] = MEM[2090] + MEM[2452];
assign MEM[2796] = MEM[2094] + MEM[1718];
assign MEM[2797] = MEM[2095] + MEM[2623];
assign MEM[2798] = MEM[2098] + MEM[2538];
assign MEM[2799] = MEM[2099] + MEM[2672];
assign MEM[2800] = MEM[2104] + MEM[2572];
assign MEM[2801] = MEM[2123] + MEM[2288];
assign MEM[2802] = MEM[2124] + MEM[2454];
assign MEM[2803] = MEM[2125] + MEM[2442];
assign MEM[2804] = MEM[2127] + MEM[2303];
assign MEM[2805] = MEM[2129] + MEM[2581];
assign MEM[2806] = MEM[2132] + MEM[2458];
assign MEM[2807] = MEM[2139] + MEM[2282];
assign MEM[2808] = MEM[2143] + MEM[2418];
assign MEM[2809] = MEM[2144] + MEM[1444];
assign MEM[2810] = MEM[2145] + MEM[2460];
assign MEM[2811] = MEM[2168] + MEM[2721];
assign MEM[2812] = MEM[2170] + MEM[1376];
assign MEM[2813] = MEM[2177] + MEM[2703];
assign MEM[2814] = MEM[2180] + MEM[2563];
assign MEM[2815] = MEM[2181] + MEM[1803];
assign MEM[2816] = MEM[2185] + MEM[1644];
assign MEM[2817] = MEM[2194] + MEM[2406];
assign MEM[2818] = MEM[2200] + MEM[2428];
assign MEM[2819] = MEM[2201] + MEM[2364];
assign MEM[2820] = MEM[2203] + MEM[2425];
assign MEM[2821] = MEM[2212] + MEM[2706];
assign MEM[2822] = MEM[2213] + MEM[2453];
assign MEM[2823] = MEM[2218] + MEM[2397];
assign MEM[2824] = MEM[2223] + MEM[1635];
assign MEM[2825] = MEM[2224] + MEM[1480];
assign MEM[2826] = MEM[2226] + MEM[1704];
assign MEM[2827] = MEM[2228] + MEM[2604];
assign MEM[2828] = MEM[2233] + MEM[2383];
assign MEM[2829] = MEM[2242] + MEM[1534];
assign MEM[2830] = MEM[2250] + MEM[2417];
assign MEM[2831] = MEM[2253] + MEM[1598];
assign MEM[2832] = MEM[2255] + MEM[1780];
assign MEM[2833] = MEM[2259] + MEM[1627];
assign MEM[2834] = MEM[2260] + MEM[1735];
assign MEM[2835] = MEM[2263] + MEM[2647];
assign MEM[2836] = MEM[2264] + MEM[2729];
assign MEM[2837] = MEM[2265] + MEM[1546];
assign MEM[2838] = MEM[2269] + MEM[2426];
assign MEM[2839] = MEM[2289] + MEM[1702];
assign MEM[2840] = MEM[2294] + MEM[2502];
assign MEM[2841] = MEM[2295] + MEM[1549];
assign MEM[2842] = MEM[2299] + MEM[2577];
assign MEM[2843] = MEM[2300] + MEM[1593];
assign MEM[2844] = MEM[2302] + MEM[1463];
assign MEM[2845] = MEM[2312] + MEM[2474];
assign MEM[2846] = MEM[2324] + MEM[2605];
assign MEM[2847] = MEM[2329] + MEM[1606];
assign MEM[2848] = MEM[2334] + MEM[1510];
assign MEM[2849] = MEM[2337] + MEM[2600];
assign MEM[2850] = MEM[2338] + MEM[1406];
assign MEM[2851] = MEM[2345] + MEM[1776];
assign MEM[2852] = MEM[2346] + MEM[2608];
assign MEM[2853] = MEM[2352] + MEM[1445];
assign MEM[2854] = MEM[2365] + MEM[1791];
assign MEM[2855] = MEM[2367] + MEM[1432];
assign MEM[2856] = MEM[2373] + MEM[2552];
assign MEM[2857] = MEM[2381] + MEM[1806];
assign MEM[2858] = MEM[2385] + MEM[2713];
assign MEM[2859] = MEM[2390] + MEM[1665];
assign MEM[2860] = MEM[2401] + MEM[2712];
assign MEM[2861] = MEM[2404] + MEM[2597];
assign MEM[2862] = MEM[2411] + MEM[2655];
assign MEM[2863] = MEM[2415] + MEM[2675];
assign MEM[2864] = MEM[2462] + MEM[2646];
assign MEM[2865] = MEM[2466] + MEM[2698];
assign MEM[2866] = MEM[2473] + MEM[1672];
assign MEM[2867] = MEM[2481] + MEM[1557];
assign MEM[2868] = MEM[2486] + MEM[2662];
assign MEM[2869] = MEM[2490] + MEM[2621];
assign MEM[2870] = MEM[2499] + MEM[1777];
assign MEM[2871] = MEM[2503] + MEM[1637];
assign MEM[2872] = MEM[2520] + MEM[1626];
assign MEM[2873] = MEM[2524] + MEM[2671];
assign MEM[2874] = MEM[2526] + MEM[1787];
assign MEM[2875] = MEM[2528] + MEM[1622];
assign MEM[2876] = MEM[2535] + MEM[2620];
assign MEM[2877] = MEM[2558] + MEM[1790];
assign MEM[2878] = MEM[2568] + MEM[1797];
assign MEM[2879] = MEM[2578] + MEM[1781];
assign MEM[2880] = MEM[2637] + MEM[2769];
assign MEM[2881] = MEM[2641] + MEM[2819];
assign MEM[2882] = MEM[2661] + MEM[1684];
assign MEM[2883] = MEM[2667] + MEM[1807];
assign MEM[2884] = MEM[2676] + MEM[2726];
assign MEM[2885] = MEM[2696] + MEM[1809];
assign MEM[2886] = MEM[2705] + MEM[2730];
assign MEM[2887] = MEM[1] + MEM[74];
assign MEM[2888] = MEM[3] + MEM[437];
assign MEM[2889] = MEM[5] + MEM[333];
assign MEM[2890] = MEM[6] + MEM[34];
assign MEM[2891] = MEM[8] + MEM[82];
assign MEM[2892] = MEM[10] + MEM[427];
assign MEM[2893] = MEM[11] + MEM[154];
assign MEM[2894] = MEM[12] + MEM[165];
assign MEM[2895] = MEM[18] + MEM[100];
assign MEM[2896] = MEM[22] + MEM[48];
assign MEM[2897] = MEM[22] + MEM[462];
assign MEM[2898] = MEM[27] + MEM[308];
assign MEM[2899] = MEM[30] + MEM[68];
assign MEM[2900] = MEM[31] + MEM[208];
assign MEM[2901] = MEM[35] + MEM[403];
assign MEM[2902] = MEM[37] + MEM[215];
assign MEM[2903] = MEM[38] + MEM[98];
assign MEM[2904] = MEM[39] + MEM[320];
assign MEM[2905] = MEM[40] + MEM[218];
assign MEM[2906] = MEM[42] + MEM[434];
assign MEM[2907] = MEM[46] + MEM[74];
assign MEM[2908] = MEM[52] + MEM[76];
assign MEM[2909] = MEM[54] + MEM[56];
assign MEM[2910] = MEM[55] + MEM[242];
assign MEM[2911] = MEM[65] + MEM[347];
assign MEM[2912] = MEM[75] + MEM[387];
assign MEM[2913] = MEM[76] + MEM[396];
assign MEM[2914] = MEM[79] + MEM[109];
assign MEM[2915] = MEM[80] + MEM[161];
assign MEM[2916] = MEM[84] + MEM[412];
assign MEM[2917] = MEM[91] + MEM[288];
assign MEM[2918] = MEM[92] + MEM[196];
assign MEM[2919] = MEM[94] + MEM[285];
assign MEM[2920] = MEM[96] + MEM[111];
assign MEM[2921] = MEM[99] + MEM[295];
assign MEM[2922] = MEM[100] + MEM[228];
assign MEM[2923] = MEM[101] + MEM[145];
assign MEM[2924] = MEM[109] + MEM[126];
assign MEM[2925] = MEM[110] + MEM[172];
assign MEM[2926] = MEM[116] + MEM[272];
assign MEM[2927] = MEM[121] + MEM[152];
assign MEM[2928] = MEM[127] + MEM[200];
assign MEM[2929] = MEM[128] + MEM[138];
assign MEM[2930] = MEM[130] + MEM[175];
assign MEM[2931] = MEM[135] + MEM[260];
assign MEM[2932] = MEM[140] + MEM[201];
assign MEM[2933] = MEM[141] + MEM[264];
assign MEM[2934] = MEM[142] + MEM[146];
assign MEM[2935] = MEM[144] + MEM[310];
assign MEM[2936] = MEM[147] + MEM[167];
assign MEM[2937] = MEM[150] + MEM[241];
assign MEM[2938] = MEM[157] + MEM[237];
assign MEM[2939] = MEM[171] + MEM[199];
assign MEM[2940] = MEM[179] + MEM[227];
assign MEM[2941] = MEM[188] + MEM[259];
assign MEM[2942] = MEM[189] + MEM[443];
assign MEM[2943] = MEM[198] + MEM[270];
assign MEM[2944] = MEM[202] + MEM[290];
assign MEM[2945] = MEM[207] + MEM[311];
assign MEM[2946] = MEM[212] + MEM[289];
assign MEM[2947] = MEM[247] + MEM[422];
assign MEM[2948] = MEM[250] + MEM[342];
assign MEM[2949] = MEM[255] + MEM[306];
assign MEM[2950] = MEM[258] + MEM[672];
assign MEM[2951] = MEM[261] + MEM[350];
assign MEM[2952] = MEM[269] + MEM[366];
assign MEM[2953] = MEM[271] + MEM[293];
assign MEM[2954] = MEM[273] + MEM[331];
assign MEM[2955] = MEM[274] + MEM[366];
assign MEM[2956] = MEM[276] + MEM[287];
assign MEM[2957] = MEM[277] + MEM[381];
assign MEM[2958] = MEM[291] + MEM[368];
assign MEM[2959] = MEM[294] + MEM[508];
assign MEM[2960] = MEM[296] + MEM[307];
assign MEM[2961] = MEM[301] + MEM[392];
assign MEM[2962] = MEM[302] + MEM[315];
assign MEM[2963] = MEM[317] + MEM[367];
assign MEM[2964] = MEM[323] + MEM[385];
assign MEM[2965] = MEM[325] + MEM[402];
assign MEM[2966] = MEM[326] + MEM[560];
assign MEM[2967] = MEM[327] + MEM[348];
assign MEM[2968] = MEM[327] + MEM[572];
assign MEM[2969] = MEM[335] + MEM[417];
assign MEM[2970] = MEM[338] + MEM[339];
assign MEM[2971] = MEM[340] + MEM[751];
assign MEM[2972] = MEM[343] + MEM[523];
assign MEM[2973] = MEM[344] + MEM[423];
assign MEM[2974] = MEM[348] + MEM[355];
assign MEM[2975] = MEM[349] + MEM[365];
assign MEM[2976] = MEM[349] + MEM[508];
assign MEM[2977] = MEM[351] + MEM[445];
assign MEM[2978] = MEM[356] + MEM[402];
assign MEM[2979] = MEM[364] + MEM[574];
assign MEM[2980] = MEM[372] + MEM[373];
assign MEM[2981] = MEM[375] + MEM[579];
assign MEM[2982] = MEM[382] + MEM[470];
assign MEM[2983] = MEM[388] + MEM[506];
assign MEM[2984] = MEM[391] + MEM[460];
assign MEM[2985] = MEM[395] + MEM[583];
assign MEM[2986] = MEM[400] + MEM[469];
assign MEM[2987] = MEM[406] + MEM[711];
assign MEM[2988] = MEM[408] + MEM[527];
assign MEM[2989] = MEM[411] + MEM[468];
assign MEM[2990] = MEM[411] + MEM[516];
assign MEM[2991] = MEM[413] + MEM[502];
assign MEM[2992] = MEM[415] + MEM[424];
assign MEM[2993] = MEM[419] + MEM[449];
assign MEM[2994] = MEM[431] + MEM[441];
assign MEM[2995] = MEM[442] + MEM[459];
assign MEM[2996] = MEM[444] + MEM[1173];
assign MEM[2997] = MEM[452] + MEM[486];
assign MEM[2998] = MEM[455] + MEM[509];
assign MEM[2999] = MEM[459] + MEM[633];
assign MEM[3000] = MEM[463] + MEM[626];
assign MEM[3001] = MEM[465] + MEM[481];
assign MEM[3002] = MEM[465] + MEM[526];
assign MEM[3003] = MEM[472] + MEM[602];
assign MEM[3004] = MEM[474] + MEM[475];
assign MEM[3005] = MEM[475] + MEM[478];
assign MEM[3006] = MEM[476] + MEM[477];
assign MEM[3007] = MEM[482] + MEM[513];
assign MEM[3008] = MEM[484] + MEM[567];
assign MEM[3009] = MEM[487] + MEM[585];
assign MEM[3010] = MEM[490] + MEM[494];
assign MEM[3011] = MEM[491] + MEM[592];
assign MEM[3012] = MEM[492] + MEM[599];
assign MEM[3013] = MEM[492] + MEM[619];
assign MEM[3014] = MEM[502] + MEM[979];
assign MEM[3015] = MEM[504] + MEM[728];
assign MEM[3016] = MEM[507] + MEM[598];
assign MEM[3017] = MEM[511] + MEM[805];
assign MEM[3018] = MEM[514] + MEM[555];
assign MEM[3019] = MEM[523] + MEM[588];
assign MEM[3020] = MEM[527] + MEM[618];
assign MEM[3021] = MEM[529] + MEM[549];
assign MEM[3022] = MEM[532] + MEM[644];
assign MEM[3023] = MEM[534] + MEM[653];
assign MEM[3024] = MEM[536] + MEM[603];
assign MEM[3025] = MEM[539] + MEM[920];
assign MEM[3026] = MEM[541] + MEM[766];
assign MEM[3027] = MEM[542] + MEM[872];
assign MEM[3028] = MEM[545] + MEM[561];
assign MEM[3029] = MEM[547] + MEM[558];
assign MEM[3030] = MEM[550] + MEM[559];
assign MEM[3031] = MEM[554] + MEM[710];
assign MEM[3032] = MEM[556] + MEM[680];
assign MEM[3033] = MEM[557] + MEM[610];
assign MEM[3034] = MEM[561] + MEM[628];
assign MEM[3035] = MEM[563] + MEM[730];
assign MEM[3036] = MEM[565] + MEM[701];
assign MEM[3037] = MEM[568] + MEM[580];
assign MEM[3038] = MEM[569] + MEM[736];
assign MEM[3039] = MEM[578] + MEM[675];
assign MEM[3040] = MEM[581] + MEM[700];
assign MEM[3041] = MEM[582] + MEM[640];
assign MEM[3042] = MEM[584] + MEM[651];
assign MEM[3043] = MEM[586] + MEM[776];
assign MEM[3044] = MEM[587] + MEM[593];
assign MEM[3045] = MEM[590] + MEM[608];
assign MEM[3046] = MEM[590] + MEM[670];
assign MEM[3047] = MEM[594] + MEM[896];
assign MEM[3048] = MEM[598] + MEM[921];
assign MEM[3049] = MEM[604] + MEM[715];
assign MEM[3050] = MEM[605] + MEM[889];
assign MEM[3051] = MEM[612] + MEM[767];
assign MEM[3052] = MEM[615] + MEM[635];
assign MEM[3053] = MEM[621] + MEM[717];
assign MEM[3054] = MEM[622] + MEM[829];
assign MEM[3055] = MEM[623] + MEM[625];
assign MEM[3056] = MEM[624] + MEM[699];
assign MEM[3057] = MEM[629] + MEM[668];
assign MEM[3058] = MEM[634] + MEM[679];
assign MEM[3059] = MEM[635] + MEM[739];
assign MEM[3060] = MEM[641] + MEM[739];
assign MEM[3061] = MEM[646] + MEM[730];
assign MEM[3062] = MEM[656] + MEM[833];
assign MEM[3063] = MEM[658] + MEM[663];
assign MEM[3064] = MEM[664] + MEM[667];
assign MEM[3065] = MEM[665] + MEM[686];
assign MEM[3066] = MEM[671] + MEM[694];
assign MEM[3067] = MEM[683] + MEM[749];
assign MEM[3068] = MEM[689] + MEM[729];
assign MEM[3069] = MEM[690] + MEM[732];
assign MEM[3070] = MEM[691] + MEM[717];
assign MEM[3071] = MEM[695] + MEM[707];
assign MEM[3072] = MEM[696] + MEM[824];
assign MEM[3073] = MEM[698] + MEM[849];
assign MEM[3074] = MEM[705] + MEM[707];
assign MEM[3075] = MEM[716] + MEM[1196];
assign MEM[3076] = MEM[718] + MEM[904];
assign MEM[3077] = MEM[734] + MEM[841];
assign MEM[3078] = MEM[735] + MEM[750];
assign MEM[3079] = MEM[740] + MEM[773];
assign MEM[3080] = MEM[741] + MEM[919];
assign MEM[3081] = MEM[744] + MEM[816];
assign MEM[3082] = MEM[747] + MEM[831];
assign MEM[3083] = MEM[750] + MEM[855];
assign MEM[3084] = MEM[751] + MEM[864];
assign MEM[3085] = MEM[752] + MEM[913];
assign MEM[3086] = MEM[753] + MEM[837];
assign MEM[3087] = MEM[754] + MEM[922];
assign MEM[3088] = MEM[755] + MEM[862];
assign MEM[3089] = MEM[756] + MEM[825];
assign MEM[3090] = MEM[757] + MEM[910];
assign MEM[3091] = MEM[760] + MEM[957];
assign MEM[3092] = MEM[765] + MEM[797];
assign MEM[3093] = MEM[767] + MEM[871];
assign MEM[3094] = MEM[770] + MEM[908];
assign MEM[3095] = MEM[770] + MEM[1009];
assign MEM[3096] = MEM[775] + MEM[788];
assign MEM[3097] = MEM[776] + MEM[842];
assign MEM[3098] = MEM[781] + MEM[823];
assign MEM[3099] = MEM[784] + MEM[1343];
assign MEM[3100] = MEM[795] + MEM[817];
assign MEM[3101] = MEM[795] + MEM[822];
assign MEM[3102] = MEM[798] + MEM[884];
assign MEM[3103] = MEM[801] + MEM[912];
assign MEM[3104] = MEM[807] + MEM[887];
assign MEM[3105] = MEM[809] + MEM[958];
assign MEM[3106] = MEM[813] + MEM[848];
assign MEM[3107] = MEM[815] + MEM[827];
assign MEM[3108] = MEM[816] + MEM[1072];
assign MEM[3109] = MEM[820] + MEM[957];
assign MEM[3110] = MEM[821] + MEM[926];
assign MEM[3111] = MEM[831] + MEM[843];
assign MEM[3112] = MEM[832] + MEM[920];
assign MEM[3113] = MEM[835] + MEM[858];
assign MEM[3114] = MEM[836] + MEM[890];
assign MEM[3115] = MEM[850] + MEM[911];
assign MEM[3116] = MEM[851] + MEM[965];
assign MEM[3117] = MEM[859] + MEM[943];
assign MEM[3118] = MEM[862] + MEM[863];
assign MEM[3119] = MEM[865] + MEM[1359];
assign MEM[3120] = MEM[868] + MEM[946];
assign MEM[3121] = MEM[869] + MEM[982];
assign MEM[3122] = MEM[870] + MEM[982];
assign MEM[3123] = MEM[875] + MEM[964];
assign MEM[3124] = MEM[876] + MEM[967];
assign MEM[3125] = MEM[878] + MEM[901];
assign MEM[3126] = MEM[878] + MEM[929];
assign MEM[3127] = MEM[881] + MEM[930];
assign MEM[3128] = MEM[882] + MEM[980];
assign MEM[3129] = MEM[884] + MEM[968];
assign MEM[3130] = MEM[889] + MEM[895];
assign MEM[3131] = MEM[893] + MEM[1223];
assign MEM[3132] = MEM[899] + MEM[941];
assign MEM[3133] = MEM[901] + MEM[951];
assign MEM[3134] = MEM[904] + MEM[1158];
assign MEM[3135] = MEM[905] + MEM[988];
assign MEM[3136] = MEM[910] + MEM[913];
assign MEM[3137] = MEM[927] + MEM[993];
assign MEM[3138] = MEM[930] + MEM[1088];
assign MEM[3139] = MEM[932] + MEM[995];
assign MEM[3140] = MEM[933] + MEM[1033];
assign MEM[3141] = MEM[937] + MEM[1053];
assign MEM[3142] = MEM[938] + MEM[975];
assign MEM[3143] = MEM[939] + MEM[998];
assign MEM[3144] = MEM[941] + MEM[956];
assign MEM[3145] = MEM[943] + MEM[966];
assign MEM[3146] = MEM[946] + MEM[1048];
assign MEM[3147] = MEM[948] + MEM[983];
assign MEM[3148] = MEM[949] + MEM[1003];
assign MEM[3149] = MEM[955] + MEM[973];
assign MEM[3150] = MEM[958] + MEM[1000];
assign MEM[3151] = MEM[960] + MEM[1066];
assign MEM[3152] = MEM[961] + MEM[981];
assign MEM[3153] = MEM[962] + MEM[985];
assign MEM[3154] = MEM[963] + MEM[1030];
assign MEM[3155] = MEM[969] + MEM[1034];
assign MEM[3156] = MEM[971] + MEM[1032];
assign MEM[3157] = MEM[976] + MEM[1061];
assign MEM[3158] = MEM[977] + MEM[1208];
assign MEM[3159] = MEM[978] + MEM[1059];
assign MEM[3160] = MEM[986] + MEM[1046];
assign MEM[3161] = MEM[986] + MEM[1071];
assign MEM[3162] = MEM[986] + MEM[1098];
assign MEM[3163] = MEM[990] + MEM[1052];
assign MEM[3164] = MEM[992] + MEM[1091];
assign MEM[3165] = MEM[993] + MEM[1039];
assign MEM[3166] = MEM[994] + MEM[1054];
assign MEM[3167] = MEM[996] + MEM[1065];
assign MEM[3168] = MEM[997] + MEM[999];
assign MEM[3169] = MEM[998] + MEM[1001];
assign MEM[3170] = MEM[998] + MEM[1296];
assign MEM[3171] = MEM[1005] + MEM[1187];
assign MEM[3172] = MEM[1007] + MEM[1008];
assign MEM[3173] = MEM[1008] + MEM[1211];
assign MEM[3174] = MEM[1011] + MEM[1024];
assign MEM[3175] = MEM[1013] + MEM[1016];
assign MEM[3176] = MEM[1015] + MEM[1038];
assign MEM[3177] = MEM[1019] + MEM[1206];
assign MEM[3178] = MEM[1021] + MEM[1162];
assign MEM[3179] = MEM[1022] + MEM[1055];
assign MEM[3180] = MEM[1025] + MEM[1036];
assign MEM[3181] = MEM[1026] + MEM[1031];
assign MEM[3182] = MEM[1030] + MEM[1068];
assign MEM[3183] = MEM[1035] + MEM[1169];
assign MEM[3184] = MEM[1037] + MEM[1141];
assign MEM[3185] = MEM[1040] + MEM[1051];
assign MEM[3186] = MEM[1042] + MEM[1043];
assign MEM[3187] = MEM[1044] + MEM[1398];
assign MEM[3188] = MEM[1045] + MEM[1066];
assign MEM[3189] = MEM[1047] + MEM[1165];
assign MEM[3190] = MEM[1049] + MEM[1127];
assign MEM[3191] = MEM[1050] + MEM[1177];
assign MEM[3192] = MEM[1052] + MEM[1147];
assign MEM[3193] = MEM[1053] + MEM[1060];
assign MEM[3194] = MEM[1053] + MEM[1193];
assign MEM[3195] = MEM[1054] + MEM[1067];
assign MEM[3196] = MEM[1054] + MEM[1225];
assign MEM[3197] = MEM[1056] + MEM[1063];
assign MEM[3198] = MEM[1057] + MEM[1129];
assign MEM[3199] = MEM[1071] + MEM[1126];
assign MEM[3200] = MEM[1074] + MEM[1130];
assign MEM[3201] = MEM[1079] + MEM[1349];
assign MEM[3202] = MEM[1080] + MEM[1089];
assign MEM[3203] = MEM[1081] + MEM[1119];
assign MEM[3204] = MEM[1082] + MEM[1110];
assign MEM[3205] = MEM[1083] + MEM[1109];
assign MEM[3206] = MEM[1085] + MEM[1183];
assign MEM[3207] = MEM[1094] + MEM[1251];
assign MEM[3208] = MEM[1095] + MEM[1152];
assign MEM[3209] = MEM[1096] + MEM[1229];
assign MEM[3210] = MEM[1099] + MEM[1148];
assign MEM[3211] = MEM[1100] + MEM[1133];
assign MEM[3212] = MEM[1101] + MEM[1216];
assign MEM[3213] = MEM[1102] + MEM[1245];
assign MEM[3214] = MEM[1103] + MEM[1427];
assign MEM[3215] = MEM[1106] + MEM[1134];
assign MEM[3216] = MEM[1115] + MEM[1118];
assign MEM[3217] = MEM[1120] + MEM[1121];
assign MEM[3218] = MEM[1122] + MEM[1123];
assign MEM[3219] = MEM[1122] + MEM[1172];
assign MEM[3220] = MEM[1135] + MEM[1137];
assign MEM[3221] = MEM[1143] + MEM[1288];
assign MEM[3222] = MEM[1144] + MEM[1157];
assign MEM[3223] = MEM[1146] + MEM[1370];
assign MEM[3224] = MEM[1154] + MEM[1245];
assign MEM[3225] = MEM[1155] + MEM[1189];
assign MEM[3226] = MEM[1155] + MEM[1668];
assign MEM[3227] = MEM[1163] + MEM[1241];
assign MEM[3228] = MEM[1167] + MEM[1193];
assign MEM[3229] = MEM[1170] + MEM[1179];
assign MEM[3230] = MEM[1170] + MEM[1192];
assign MEM[3231] = MEM[1170] + MEM[1215];
assign MEM[3232] = MEM[1173] + MEM[1242];
assign MEM[3233] = MEM[1173] + MEM[1283];
assign MEM[3234] = MEM[1175] + MEM[1381];
assign MEM[3235] = MEM[1181] + MEM[1251];
assign MEM[3236] = MEM[1182] + MEM[1197];
assign MEM[3237] = MEM[1183] + MEM[1365];
assign MEM[3238] = MEM[1183] + MEM[1378];
assign MEM[3239] = MEM[1184] + MEM[1229];
assign MEM[3240] = MEM[1185] + MEM[1186];
assign MEM[3241] = MEM[1186] + MEM[1199];
assign MEM[3242] = MEM[1186] + MEM[1202];
assign MEM[3243] = MEM[1188] + MEM[1212];
assign MEM[3244] = MEM[1192] + MEM[1317];
assign MEM[3245] = MEM[1192] + MEM[1404];
assign MEM[3246] = MEM[1195] + MEM[1209];
assign MEM[3247] = MEM[1200] + MEM[1203];
assign MEM[3248] = MEM[1203] + MEM[1230];
assign MEM[3249] = MEM[1204] + MEM[1249];
assign MEM[3250] = MEM[1205] + MEM[1342];
assign MEM[3251] = MEM[1207] + MEM[1318];
assign MEM[3252] = MEM[1210] + MEM[1219];
assign MEM[3253] = MEM[1213] + MEM[1277];
assign MEM[3254] = MEM[1214] + MEM[1272];
assign MEM[3255] = MEM[1217] + MEM[1267];
assign MEM[3256] = MEM[1218] + MEM[1359];
assign MEM[3257] = MEM[1222] + MEM[1228];
assign MEM[3258] = MEM[1228] + MEM[1260];
assign MEM[3259] = MEM[1237] + MEM[1346];
assign MEM[3260] = MEM[1241] + MEM[1242];
assign MEM[3261] = MEM[1249] + MEM[1441];
assign MEM[3262] = MEM[1255] + MEM[1300];
assign MEM[3263] = MEM[1260] + MEM[1470];
assign MEM[3264] = MEM[1263] + MEM[1270];
assign MEM[3265] = MEM[1263] + MEM[1407];
assign MEM[3266] = MEM[1265] + MEM[1377];
assign MEM[3267] = MEM[1265] + MEM[1422];
assign MEM[3268] = MEM[1267] + MEM[1316];
assign MEM[3269] = MEM[1269] + MEM[1277];
assign MEM[3270] = MEM[1269] + MEM[1301];
assign MEM[3271] = MEM[1270] + MEM[1379];
assign MEM[3272] = MEM[1272] + MEM[1394];
assign MEM[3273] = MEM[1283] + MEM[1368];
assign MEM[3274] = MEM[1286] + MEM[1365];
assign MEM[3275] = MEM[1286] + MEM[1393];
assign MEM[3276] = MEM[1288] + MEM[1407];
assign MEM[3277] = MEM[1291] + MEM[1308];
assign MEM[3278] = MEM[1291] + MEM[1337];
assign MEM[3279] = MEM[1296] + MEM[1342];
assign MEM[3280] = MEM[1298] + MEM[1411];
assign MEM[3281] = MEM[1301] + MEM[1361];
assign MEM[3282] = MEM[1308] + MEM[1324];
assign MEM[3283] = MEM[1316] + MEM[1324];
assign MEM[3284] = MEM[1317] + MEM[1426];
assign MEM[3285] = MEM[1318] + MEM[1405];
assign MEM[3286] = MEM[1331] + MEM[1358];
assign MEM[3287] = MEM[1331] + MEM[1384];
assign MEM[3288] = MEM[1337] + MEM[1348];
assign MEM[3289] = MEM[1343] + MEM[1400];
assign MEM[3290] = MEM[1346] + MEM[1350];
assign MEM[3291] = MEM[1348] + MEM[1475];
assign MEM[3292] = MEM[1349] + MEM[1421];
assign MEM[3293] = MEM[1350] + MEM[1450];
assign MEM[3294] = MEM[1358] + MEM[1502];
assign MEM[3295] = MEM[1361] + MEM[1415];
assign MEM[3296] = MEM[1366] + MEM[1390];
assign MEM[3297] = MEM[1366] + MEM[1409];
assign MEM[3298] = MEM[1367] + MEM[1399];
assign MEM[3299] = MEM[1367] + MEM[1425];
assign MEM[3300] = MEM[1368] + MEM[1477];
assign MEM[3301] = MEM[1370] + MEM[1442];
assign MEM[3302] = MEM[1376] + MEM[1431];
assign MEM[3303] = MEM[1380] + MEM[1476];
assign MEM[3304] = MEM[1382] + MEM[1407];
assign MEM[3305] = MEM[1383] + MEM[1453];
assign MEM[3306] = MEM[1385] + MEM[1494];
assign MEM[3307] = MEM[1387] + MEM[1452];
assign MEM[3308] = MEM[1388] + MEM[1409];
assign MEM[3309] = MEM[1389] + MEM[1409];
assign MEM[3310] = MEM[1391] + MEM[1446];
assign MEM[3311] = MEM[1392] + MEM[1401];
assign MEM[3312] = MEM[1395] + MEM[1412];
assign MEM[3313] = MEM[1396] + MEM[1455];
assign MEM[3314] = MEM[1397] + MEM[1424];
assign MEM[3315] = MEM[1402] + MEM[1434];
assign MEM[3316] = MEM[1403] + MEM[1451];
assign MEM[3317] = MEM[1406] + MEM[1457];
assign MEM[3318] = MEM[1408] + MEM[1480];
assign MEM[3319] = MEM[1410] + MEM[1539];
assign MEM[3320] = MEM[1412] + MEM[1416];
assign MEM[3321] = MEM[1412] + MEM[1533];
assign MEM[3322] = MEM[1413] + MEM[1526];
assign MEM[3323] = MEM[1414] + MEM[1461];
assign MEM[3324] = MEM[1418] + MEM[1448];
assign MEM[3325] = MEM[1419] + MEM[1443];
assign MEM[3326] = MEM[1423] + MEM[1537];
assign MEM[3327] = MEM[1428] + MEM[1512];
assign MEM[3328] = MEM[1429] + MEM[1478];
assign MEM[3329] = MEM[1430] + MEM[1482];
assign MEM[3330] = MEM[1431] + MEM[1459];
assign MEM[3331] = MEM[1431] + MEM[1573];
assign MEM[3332] = MEM[1432] + MEM[1513];
assign MEM[3333] = MEM[1433] + MEM[1463];
assign MEM[3334] = MEM[1435] + MEM[1467];
assign MEM[3335] = MEM[1436] + MEM[1554];
assign MEM[3336] = MEM[1437] + MEM[1442];
assign MEM[3337] = MEM[1438] + MEM[1517];
assign MEM[3338] = MEM[1439] + MEM[1524];
assign MEM[3339] = MEM[1440] + MEM[1465];
assign MEM[3340] = MEM[1441] + MEM[1492];
assign MEM[3341] = MEM[1441] + MEM[1570];
assign MEM[3342] = MEM[1442] + MEM[1737];
assign MEM[3343] = MEM[1444] + MEM[1550];
assign MEM[3344] = MEM[1445] + MEM[1633];
assign MEM[3345] = MEM[1447] + MEM[1490];
assign MEM[3346] = MEM[1449] + MEM[1505];
assign MEM[3347] = MEM[1454] + MEM[1490];
assign MEM[3348] = MEM[1456] + MEM[1486];
assign MEM[3349] = MEM[1458] + MEM[1464];
assign MEM[3350] = MEM[1460] + MEM[1479];
assign MEM[3351] = MEM[1468] + MEM[1549];
assign MEM[3352] = MEM[1469] + MEM[1496];
assign MEM[3353] = MEM[1471] + MEM[1590];
assign MEM[3354] = MEM[1472] + MEM[1571];
assign MEM[3355] = MEM[1473] + MEM[1628];
assign MEM[3356] = MEM[1474] + MEM[1519];
assign MEM[3357] = MEM[1476] + MEM[1495];
assign MEM[3358] = MEM[1476] + MEM[1548];
assign MEM[3359] = MEM[1479] + MEM[1538];
assign MEM[3360] = MEM[1479] + MEM[1560];
assign MEM[3361] = MEM[1481] + MEM[1553];
assign MEM[3362] = MEM[1483] + MEM[1490];
assign MEM[3363] = MEM[1484] + MEM[1539];
assign MEM[3364] = MEM[1485] + MEM[1532];
assign MEM[3365] = MEM[1487] + MEM[1659];
assign MEM[3366] = MEM[1488] + MEM[1558];
assign MEM[3367] = MEM[1489] + MEM[1493];
assign MEM[3368] = MEM[1491] + MEM[1547];
assign MEM[3369] = MEM[1493] + MEM[1552];
assign MEM[3370] = MEM[1493] + MEM[1605];
assign MEM[3371] = MEM[1497] + MEM[1522];
assign MEM[3372] = MEM[1498] + MEM[1694];
assign MEM[3373] = MEM[1499] + MEM[1569];
assign MEM[3374] = MEM[1500] + MEM[1534];
assign MEM[3375] = MEM[1504] + MEM[1636];
assign MEM[3376] = MEM[1506] + MEM[1784];
assign MEM[3377] = MEM[1507] + MEM[1567];
assign MEM[3378] = MEM[1508] + MEM[1650];
assign MEM[3379] = MEM[1509] + MEM[1656];
assign MEM[3380] = MEM[1510] + MEM[1579];
assign MEM[3381] = MEM[1511] + MEM[1609];
assign MEM[3382] = MEM[1514] + MEM[1525];
assign MEM[3383] = MEM[1515] + MEM[1816];
assign MEM[3384] = MEM[1516] + MEM[1592];
assign MEM[3385] = MEM[1518] + MEM[1578];
assign MEM[3386] = MEM[1520] + MEM[1755];
assign MEM[3387] = MEM[1521] + MEM[1652];
assign MEM[3388] = MEM[1523] + MEM[1567];
assign MEM[3389] = MEM[1527] + MEM[1721];
assign MEM[3390] = MEM[1528] + MEM[1535];
assign MEM[3391] = MEM[1529] + MEM[1581];
assign MEM[3392] = MEM[1530] + MEM[1628];
assign MEM[3393] = MEM[1531] + MEM[1541];
assign MEM[3394] = MEM[1533] + MEM[1555];
assign MEM[3395] = MEM[1533] + MEM[1577];
assign MEM[3396] = MEM[1536] + MEM[1611];
assign MEM[3397] = MEM[1539] + MEM[1597];
assign MEM[3398] = MEM[1540] + MEM[1562];
assign MEM[3399] = MEM[1542] + MEM[1623];
assign MEM[3400] = MEM[1543] + MEM[1557];
assign MEM[3401] = MEM[1544] + MEM[1651];
assign MEM[3402] = MEM[1545] + MEM[1632];
assign MEM[3403] = MEM[1546] + MEM[1608];
assign MEM[3404] = MEM[1551] + MEM[1572];
assign MEM[3405] = MEM[1556] + MEM[1576];
assign MEM[3406] = MEM[1561] + MEM[1663];
assign MEM[3407] = MEM[1563] + MEM[1624];
assign MEM[3408] = MEM[1564] + MEM[1589];
assign MEM[3409] = MEM[1565] + MEM[1647];
assign MEM[3410] = MEM[1566] + MEM[1595];
assign MEM[3411] = MEM[1567] + MEM[1604];
assign MEM[3412] = MEM[1574] + MEM[1640];
assign MEM[3413] = MEM[1575] + MEM[1724];
assign MEM[3414] = MEM[1577] + MEM[1645];
assign MEM[3415] = MEM[1577] + MEM[1813];
assign MEM[3416] = MEM[1580] + MEM[1594];
assign MEM[3417] = MEM[1582] + MEM[1684];
assign MEM[3418] = MEM[1583] + MEM[1669];
assign MEM[3419] = MEM[1584] + MEM[1588];
assign MEM[3420] = MEM[1585] + MEM[1671];
assign MEM[3421] = MEM[1586] + MEM[1662];
assign MEM[3422] = MEM[1587] + MEM[1615];
assign MEM[3423] = MEM[1591] + MEM[1676];
assign MEM[3424] = MEM[1593] + MEM[1613];
assign MEM[3425] = MEM[1595] + MEM[1602];
assign MEM[3426] = MEM[1595] + MEM[1658];
assign MEM[3427] = MEM[1596] + MEM[1613];
assign MEM[3428] = MEM[1598] + MEM[1617];
assign MEM[3429] = MEM[1599] + MEM[1635];
assign MEM[3430] = MEM[1600] + MEM[1827];
assign MEM[3431] = MEM[1601] + MEM[1770];
assign MEM[3432] = MEM[1603] + MEM[1638];
assign MEM[3433] = MEM[1606] + MEM[1622];
assign MEM[3434] = MEM[1607] + MEM[1620];
assign MEM[3435] = MEM[1609] + MEM[1678];
assign MEM[3436] = MEM[1609] + MEM[1760];
assign MEM[3437] = MEM[1610] + MEM[1671];
assign MEM[3438] = MEM[1612] + MEM[1847];
assign MEM[3439] = MEM[1613] + MEM[1619];
assign MEM[3440] = MEM[1614] + MEM[1711];
assign MEM[3441] = MEM[1616] + MEM[1628];
assign MEM[3442] = MEM[1617] + MEM[1626];
assign MEM[3443] = MEM[1617] + MEM[1706];
assign MEM[3444] = MEM[1618] + MEM[1701];
assign MEM[3445] = MEM[1621] + MEM[1657];
assign MEM[3446] = MEM[1627] + MEM[1706];
assign MEM[3447] = MEM[1629] + MEM[1689];
assign MEM[3448] = MEM[1630] + MEM[1663];
assign MEM[3449] = MEM[1631] + MEM[1739];
assign MEM[3450] = MEM[1634] + MEM[1643];
assign MEM[3451] = MEM[1637] + MEM[1706];
assign MEM[3452] = MEM[1641] + MEM[1646];
assign MEM[3453] = MEM[1642] + MEM[1661];
assign MEM[3454] = MEM[1644] + MEM[1690];
assign MEM[3455] = MEM[1648] + MEM[1817];
assign MEM[3456] = MEM[1649] + MEM[1717];
assign MEM[3457] = MEM[1653] + MEM[1696];
assign MEM[3458] = MEM[1654] + MEM[1665];
assign MEM[3459] = MEM[1655] + MEM[1674];
assign MEM[3460] = MEM[1660] + MEM[1745];
assign MEM[3461] = MEM[1663] + MEM[1757];
assign MEM[3462] = MEM[1666] + MEM[1727];
assign MEM[3463] = MEM[1667] + MEM[1672];
assign MEM[3464] = MEM[1667] + MEM[1728];
assign MEM[3465] = MEM[1667] + MEM[1730];
assign MEM[3466] = MEM[1670] + MEM[1729];
assign MEM[3467] = MEM[1671] + MEM[1780];
assign MEM[3468] = MEM[1673] + MEM[1890];
assign MEM[3469] = MEM[1674] + MEM[1699];
assign MEM[3470] = MEM[1674] + MEM[1726];
assign MEM[3471] = MEM[1675] + MEM[1770];
assign MEM[3472] = MEM[1677] + MEM[1769];
assign MEM[3473] = MEM[1679] + MEM[1802];
assign MEM[3474] = MEM[1681] + MEM[1948];
assign MEM[3475] = MEM[1682] + MEM[1897];
assign MEM[3476] = MEM[1683] + MEM[1716];
assign MEM[3477] = MEM[1685] + MEM[1846];
assign MEM[3478] = MEM[1687] + MEM[1809];
assign MEM[3479] = MEM[1688] + MEM[1723];
assign MEM[3480] = MEM[1691] + MEM[1740];
assign MEM[3481] = MEM[1692] + MEM[1719];
assign MEM[3482] = MEM[1693] + MEM[1710];
assign MEM[3483] = MEM[1695] + MEM[1699];
assign MEM[3484] = MEM[1697] + MEM[1814];
assign MEM[3485] = MEM[1698] + MEM[1709];
assign MEM[3486] = MEM[1699] + MEM[1757];
assign MEM[3487] = MEM[1700] + MEM[1766];
assign MEM[3488] = MEM[1702] + MEM[1732];
assign MEM[3489] = MEM[1703] + MEM[1758];
assign MEM[3490] = MEM[1704] + MEM[1778];
assign MEM[3491] = MEM[1705] + MEM[1738];
assign MEM[3492] = MEM[1707] + MEM[1710];
assign MEM[3493] = MEM[1708] + MEM[1718];
assign MEM[3494] = MEM[1710] + MEM[1720];
assign MEM[3495] = MEM[1712] + MEM[1725];
assign MEM[3496] = MEM[1713] + MEM[1744];
assign MEM[3497] = MEM[1714] + MEM[1742];
assign MEM[3498] = MEM[1715] + MEM[1750];
assign MEM[3499] = MEM[1722] + MEM[1731];
assign MEM[3500] = MEM[1732] + MEM[1746];
assign MEM[3501] = MEM[1732] + MEM[1882];
assign MEM[3502] = MEM[1734] + MEM[1743];
assign MEM[3503] = MEM[1735] + MEM[1778];
assign MEM[3504] = MEM[1739] + MEM[1747];
assign MEM[3505] = MEM[1739] + MEM[1778];
assign MEM[3506] = MEM[1741] + MEM[1764];
assign MEM[3507] = MEM[1747] + MEM[1751];
assign MEM[3508] = MEM[1747] + MEM[1771];
assign MEM[3509] = MEM[1748] + MEM[1766];
assign MEM[3510] = MEM[1749] + MEM[1753];
assign MEM[3511] = MEM[1752] + MEM[1829];
assign MEM[3512] = MEM[1754] + MEM[1847];
assign MEM[3513] = MEM[1756] + MEM[1760];
assign MEM[3514] = MEM[1757] + MEM[1767];
assign MEM[3515] = MEM[1759] + MEM[1896];
assign MEM[3516] = MEM[1760] + MEM[1766];
assign MEM[3517] = MEM[1761] + MEM[1824];
assign MEM[3518] = MEM[1762] + MEM[1765];
assign MEM[3519] = MEM[1763] + MEM[1765];
assign MEM[3520] = MEM[1765] + MEM[1790];
assign MEM[3521] = MEM[1769] + MEM[1770];
assign MEM[3522] = MEM[1769] + MEM[1808];
assign MEM[3523] = MEM[1772] + MEM[1774];
assign MEM[3524] = MEM[1773] + MEM[1831];
assign MEM[3525] = MEM[1774] + MEM[1789];
assign MEM[3526] = MEM[1774] + MEM[1811];
assign MEM[3527] = MEM[1775] + MEM[1805];
assign MEM[3528] = MEM[1776] + MEM[1825];
assign MEM[3529] = MEM[1777] + MEM[1812];
assign MEM[3530] = MEM[1779] + MEM[1822];
assign MEM[3531] = MEM[1781] + MEM[1791];
assign MEM[3532] = MEM[1782] + MEM[1840];
assign MEM[3533] = MEM[1783] + MEM[1788];
assign MEM[3534] = MEM[1785] + MEM[1786];
assign MEM[3535] = MEM[1785] + MEM[1797];
assign MEM[3536] = MEM[1785] + MEM[1866];
assign MEM[3537] = MEM[1787] + MEM[1822];
assign MEM[3538] = MEM[1792] + MEM[1820];
assign MEM[3539] = MEM[1793] + MEM[1794];
assign MEM[3540] = MEM[1795] + MEM[1834];
assign MEM[3541] = MEM[1796] + MEM[1919];
assign MEM[3542] = MEM[1798] + MEM[1896];
assign MEM[3543] = MEM[1799] + MEM[1889];
assign MEM[3544] = MEM[1800] + MEM[1842];
assign MEM[3545] = MEM[1801] + MEM[1875];
assign MEM[3546] = MEM[1802] + MEM[1817];
assign MEM[3547] = MEM[1802] + MEM[1904];
assign MEM[3548] = MEM[1803] + MEM[1862];
assign MEM[3549] = MEM[1804] + MEM[1881];
assign MEM[3550] = MEM[1806] + MEM[1854];
assign MEM[3551] = MEM[1807] + MEM[1810];
assign MEM[3552] = MEM[1813] + MEM[1826];
assign MEM[3553] = MEM[1813] + MEM[1894];
assign MEM[3554] = MEM[1815] + MEM[1821];
assign MEM[3555] = MEM[1816] + MEM[1818];
assign MEM[3556] = MEM[1818] + MEM[1903];
assign MEM[3557] = MEM[1820] + MEM[1825];
assign MEM[3558] = MEM[1821] + MEM[1877];
assign MEM[3559] = MEM[1824] + MEM[1829];
assign MEM[3560] = MEM[1826] + MEM[1841];
assign MEM[3561] = MEM[1827] + MEM[1899];
assign MEM[3562] = MEM[1828] + MEM[1835];
assign MEM[3563] = MEM[1828] + MEM[1874];
assign MEM[3564] = MEM[1831] + MEM[1878];
assign MEM[3565] = MEM[1834] + MEM[1866];
assign MEM[3566] = MEM[1835] + MEM[1947];
assign MEM[3567] = MEM[1836] + MEM[1900];
assign MEM[3568] = MEM[1836] + MEM[1905];
assign MEM[3569] = MEM[1837] + MEM[1845];
assign MEM[3570] = MEM[1837] + MEM[1889];
assign MEM[3571] = MEM[1838] + MEM[1875];
assign MEM[3572] = MEM[1838] + MEM[1884];
assign MEM[3573] = MEM[1840] + MEM[1860];
assign MEM[3574] = MEM[1841] + MEM[1855];
assign MEM[3575] = MEM[1842] + MEM[1880];
assign MEM[3576] = MEM[1845] + MEM[1868];
assign MEM[3577] = MEM[1846] + MEM[1867];
assign MEM[3578] = MEM[1854] + MEM[1858];
assign MEM[3579] = MEM[1855] + MEM[1939];
assign MEM[3580] = MEM[1856] + MEM[1879];
assign MEM[3581] = MEM[1856] + MEM[1880];
assign MEM[3582] = MEM[1858] + MEM[1892];
assign MEM[3583] = MEM[1860] + MEM[1901];
assign MEM[3584] = MEM[1862] + MEM[1878];
assign MEM[3585] = MEM[1865] + MEM[1886];
assign MEM[3586] = MEM[1865] + MEM[1901];
assign MEM[3587] = MEM[1867] + MEM[1996];
assign MEM[3588] = MEM[1868] + MEM[1874];
assign MEM[3589] = MEM[1871] + MEM[1885];
assign MEM[3590] = MEM[1871] + MEM[1893];
assign MEM[3591] = MEM[1873] + MEM[1884];
assign MEM[3592] = MEM[1873] + MEM[1929];
assign MEM[3593] = MEM[1877] + MEM[2153];
assign MEM[3594] = MEM[1879] + MEM[2064];
assign MEM[3595] = MEM[1881] + MEM[2047];
assign MEM[3596] = MEM[1882] + MEM[1883];
assign MEM[3597] = MEM[1883] + MEM[1888];
assign MEM[3598] = MEM[1885] + MEM[1951];
assign MEM[3599] = MEM[1886] + MEM[1951];
assign MEM[3600] = MEM[1888] + MEM[2038];
assign MEM[3601] = MEM[1890] + MEM[1935];
assign MEM[3602] = MEM[1892] + MEM[1895];
assign MEM[3603] = MEM[1893] + MEM[1912];
assign MEM[3604] = MEM[1894] + MEM[1971];
assign MEM[3605] = MEM[1895] + MEM[1898];
assign MEM[3606] = MEM[1897] + MEM[1920];
assign MEM[3607] = MEM[1898] + MEM[1933];
assign MEM[3608] = MEM[1899] + MEM[1928];
assign MEM[3609] = MEM[1900] + MEM[1999];
assign MEM[3610] = MEM[1902] + MEM[1929];
assign MEM[3611] = MEM[1902] + MEM[1973];
assign MEM[3612] = MEM[1903] + MEM[1968];
assign MEM[3613] = MEM[1904] + MEM[1907];
assign MEM[3614] = MEM[1905] + MEM[1932];
assign MEM[3615] = MEM[1906] + MEM[1915];
assign MEM[3616] = MEM[1906] + MEM[1922];
assign MEM[3617] = MEM[1907] + MEM[1928];
assign MEM[3618] = MEM[1912] + MEM[1977];
assign MEM[3619] = MEM[1915] + MEM[2027];
assign MEM[3620] = MEM[1919] + MEM[1936];
assign MEM[3621] = MEM[1920] + MEM[1936];
assign MEM[3622] = MEM[1922] + MEM[1961];
assign MEM[3623] = MEM[1925] + MEM[1938];
assign MEM[3624] = MEM[1925] + MEM[2061];
assign MEM[3625] = MEM[1927] + MEM[1953];
assign MEM[3626] = MEM[1927] + MEM[1956];
assign MEM[3627] = MEM[1932] + MEM[1967];
assign MEM[3628] = MEM[1933] + MEM[2000];
assign MEM[3629] = MEM[1935] + MEM[1938];
assign MEM[3630] = MEM[1939] + MEM[1961];
assign MEM[3631] = MEM[1943] + MEM[1946];
assign MEM[3632] = MEM[1943] + MEM[1986];
assign MEM[3633] = MEM[1944] + MEM[1976];
assign MEM[3634] = MEM[1944] + MEM[2014];
assign MEM[3635] = MEM[1946] + MEM[2103];
assign MEM[3636] = MEM[1947] + MEM[1958];
assign MEM[3637] = MEM[1948] + MEM[2008];
assign MEM[3638] = MEM[1950] + MEM[1969];
assign MEM[3639] = MEM[1950] + MEM[1970];
assign MEM[3640] = MEM[1952] + MEM[1990];
assign MEM[3641] = MEM[1952] + MEM[2022];
assign MEM[3642] = MEM[1953] + MEM[1987];
assign MEM[3643] = MEM[1956] + MEM[2059];
assign MEM[3644] = MEM[1957] + MEM[1990];
assign MEM[3645] = MEM[1957] + MEM[2061];
assign MEM[3646] = MEM[1958] + MEM[1985];
assign MEM[3647] = MEM[1962] + MEM[1966];
assign MEM[3648] = MEM[1962] + MEM[1995];
assign MEM[3649] = MEM[1964] + MEM[1971];
assign MEM[3650] = MEM[1964] + MEM[2112];
assign MEM[3651] = MEM[1966] + MEM[2081];
assign MEM[3652] = MEM[1967] + MEM[2037];
assign MEM[3653] = MEM[1968] + MEM[1998];
assign MEM[3654] = MEM[1969] + MEM[1975];
assign MEM[3655] = MEM[1970] + MEM[2010];
assign MEM[3656] = MEM[1973] + MEM[1992];
assign MEM[3657] = MEM[1975] + MEM[1978];
assign MEM[3658] = MEM[1976] + MEM[1999];
assign MEM[3659] = MEM[1977] + MEM[1987];
assign MEM[3660] = MEM[1978] + MEM[2063];
assign MEM[3661] = MEM[1985] + MEM[1988];
assign MEM[3662] = MEM[1986] + MEM[2111];
assign MEM[3663] = MEM[1988] + MEM[2037];
assign MEM[3664] = MEM[1991] + MEM[2014];
assign MEM[3665] = MEM[1991] + MEM[2024];
assign MEM[3666] = MEM[1992] + MEM[2058];
assign MEM[3667] = MEM[1993] + MEM[2017];
assign MEM[3668] = MEM[1993] + MEM[2051];
assign MEM[3669] = MEM[1995] + MEM[2045];
assign MEM[3670] = MEM[1996] + MEM[2003];
assign MEM[3671] = MEM[1998] + MEM[2031];
assign MEM[3672] = MEM[2000] + MEM[2047];
assign MEM[3673] = MEM[2001] + MEM[2010];
assign MEM[3674] = MEM[2001] + MEM[2102];
assign MEM[3675] = MEM[2003] + MEM[2060];
assign MEM[3676] = MEM[2007] + MEM[2093];
assign MEM[3677] = MEM[2007] + MEM[2119];
assign MEM[3678] = MEM[2008] + MEM[2021];
assign MEM[3679] = MEM[2009] + MEM[2027];
assign MEM[3680] = MEM[2009] + MEM[2142];
assign MEM[3681] = MEM[2012] + MEM[2035];
assign MEM[3682] = MEM[2012] + MEM[2046];
assign MEM[3683] = MEM[2016] + MEM[2028];
assign MEM[3684] = MEM[2016] + MEM[2074];
assign MEM[3685] = MEM[2017] + MEM[2038];
assign MEM[3686] = MEM[2018] + MEM[2019];
assign MEM[3687] = MEM[2018] + MEM[2138];
assign MEM[3688] = MEM[2019] + MEM[2020];
assign MEM[3689] = MEM[2020] + MEM[2199];
assign MEM[3690] = MEM[2021] + MEM[2146];
assign MEM[3691] = MEM[2022] + MEM[2262];
assign MEM[3692] = MEM[2023] + MEM[2033];
assign MEM[3693] = MEM[2023] + MEM[2075];
assign MEM[3694] = MEM[2024] + MEM[2080];
assign MEM[3695] = MEM[2028] + MEM[2058];
assign MEM[3696] = MEM[2030] + MEM[2045];
assign MEM[3697] = MEM[2030] + MEM[2204];
assign MEM[3698] = MEM[2031] + MEM[2033];
assign MEM[3699] = MEM[2032] + MEM[2075];
assign MEM[3700] = MEM[2032] + MEM[2076];
assign MEM[3701] = MEM[2035] + MEM[2051];
assign MEM[3702] = MEM[2046] + MEM[2150];
assign MEM[3703] = MEM[2048] + MEM[2097];
assign MEM[3704] = MEM[2048] + MEM[2100];
assign MEM[3705] = MEM[2052] + MEM[2065];
assign MEM[3706] = MEM[2052] + MEM[2082];
assign MEM[3707] = MEM[2056] + MEM[2065];
assign MEM[3708] = MEM[2056] + MEM[2192];
assign MEM[3709] = MEM[2059] + MEM[2072];
assign MEM[3710] = MEM[2060] + MEM[2074];
assign MEM[3711] = MEM[2063] + MEM[2067];
assign MEM[3712] = MEM[2064] + MEM[2076];
assign MEM[3713] = MEM[2066] + MEM[2096];
assign MEM[3714] = MEM[2066] + MEM[2138];
assign MEM[3715] = MEM[2067] + MEM[2069];
assign MEM[3716] = MEM[2069] + MEM[2155];
assign MEM[3717] = MEM[2070] + MEM[2173];
assign MEM[3718] = MEM[2070] + MEM[2198];
assign MEM[3719] = MEM[2072] + MEM[2150];
assign MEM[3720] = MEM[2077] + MEM[2135];
assign MEM[3721] = MEM[2077] + MEM[2149];
assign MEM[3722] = MEM[2078] + MEM[2081];
assign MEM[3723] = MEM[2078] + MEM[2103];
assign MEM[3724] = MEM[2080] + MEM[2091];
assign MEM[3725] = MEM[2082] + MEM[2088];
assign MEM[3726] = MEM[2086] + MEM[2118];
assign MEM[3727] = MEM[2086] + MEM[2146];
assign MEM[3728] = MEM[2087] + MEM[2108];
assign MEM[3729] = MEM[2087] + MEM[2128];
assign MEM[3730] = MEM[2088] + MEM[2100];
assign MEM[3731] = MEM[2091] + MEM[2097];
assign MEM[3732] = MEM[2092] + MEM[2101];
assign MEM[3733] = MEM[2092] + MEM[2210];
assign MEM[3734] = MEM[2093] + MEM[2198];
assign MEM[3735] = MEM[2096] + MEM[2130];
assign MEM[3736] = MEM[2101] + MEM[2130];
assign MEM[3737] = MEM[2102] + MEM[2111];
assign MEM[3738] = MEM[2105] + MEM[2113];
assign MEM[3739] = MEM[2105] + MEM[2126];
assign MEM[3740] = MEM[2106] + MEM[2186];
assign MEM[3741] = MEM[2106] + MEM[2199];
assign MEM[3742] = MEM[2108] + MEM[2115];
assign MEM[3743] = MEM[2109] + MEM[2113];
assign MEM[3744] = MEM[2109] + MEM[2247];
assign MEM[3745] = MEM[2110] + MEM[2154];
assign MEM[3746] = MEM[2110] + MEM[2189];
assign MEM[3747] = MEM[2112] + MEM[2131];
assign MEM[3748] = MEM[2115] + MEM[2117];
assign MEM[3749] = MEM[2117] + MEM[2159];
assign MEM[3750] = MEM[2118] + MEM[2193];
assign MEM[3751] = MEM[2119] + MEM[2135];
assign MEM[3752] = MEM[2120] + MEM[2173];
assign MEM[3753] = MEM[2120] + MEM[2219];
assign MEM[3754] = MEM[2126] + MEM[2186];
assign MEM[3755] = MEM[2128] + MEM[2234];
assign MEM[3756] = MEM[2131] + MEM[2217];
assign MEM[3757] = MEM[2136] + MEM[2141];
assign MEM[3758] = MEM[2136] + MEM[2151];
assign MEM[3759] = MEM[2137] + MEM[2158];
assign MEM[3760] = MEM[2137] + MEM[2164];
assign MEM[3761] = MEM[2141] + MEM[2214];
assign MEM[3762] = MEM[2142] + MEM[2184];
assign MEM[3763] = MEM[2147] + MEM[2158];
assign MEM[3764] = MEM[2147] + MEM[2176];
assign MEM[3765] = MEM[2148] + MEM[2156];
assign MEM[3766] = MEM[2148] + MEM[2188];
assign MEM[3767] = MEM[2149] + MEM[2160];
assign MEM[3768] = MEM[2151] + MEM[2237];
assign MEM[3769] = MEM[2153] + MEM[2360];
assign MEM[3770] = MEM[2154] + MEM[2175];
assign MEM[3771] = MEM[2155] + MEM[2193];
assign MEM[3772] = MEM[2156] + MEM[2239];
assign MEM[3773] = MEM[2157] + MEM[2179];
assign MEM[3774] = MEM[2157] + MEM[2190];
assign MEM[3775] = MEM[2159] + MEM[2206];
assign MEM[3776] = MEM[2160] + MEM[2163];
assign MEM[3777] = MEM[2162] + MEM[2284];
assign MEM[3778] = MEM[2162] + MEM[2310];
assign MEM[3779] = MEM[2163] + MEM[2174];
assign MEM[3780] = MEM[2164] + MEM[2172];
assign MEM[3781] = MEM[2166] + MEM[2189];
assign MEM[3782] = MEM[2166] + MEM[2285];
assign MEM[3783] = MEM[2171] + MEM[2178];
assign MEM[3784] = MEM[2171] + MEM[2225];
assign MEM[3785] = MEM[2172] + MEM[2191];
assign MEM[3786] = MEM[2174] + MEM[2195];
assign MEM[3787] = MEM[2175] + MEM[2243];
assign MEM[3788] = MEM[2176] + MEM[2190];
assign MEM[3789] = MEM[2178] + MEM[2267];
assign MEM[3790] = MEM[2179] + MEM[2275];
assign MEM[3791] = MEM[2183] + MEM[2187];
assign MEM[3792] = MEM[2183] + MEM[2240];
assign MEM[3793] = MEM[2184] + MEM[2419];
assign MEM[3794] = MEM[2187] + MEM[2292];
assign MEM[3795] = MEM[2188] + MEM[2215];
assign MEM[3796] = MEM[2191] + MEM[2216];
assign MEM[3797] = MEM[2192] + MEM[2221];
assign MEM[3798] = MEM[2195] + MEM[2214];
assign MEM[3799] = MEM[2196] + MEM[2230];
assign MEM[3800] = MEM[2196] + MEM[2343];
assign MEM[3801] = MEM[2202] + MEM[2215];
assign MEM[3802] = MEM[2202] + MEM[2297];
assign MEM[3803] = MEM[2204] + MEM[2231];
assign MEM[3804] = MEM[2205] + MEM[2234];
assign MEM[3805] = MEM[2205] + MEM[2283];
assign MEM[3806] = MEM[2206] + MEM[2347];
assign MEM[3807] = MEM[2207] + MEM[2208];
assign MEM[3808] = MEM[2207] + MEM[2217];
assign MEM[3809] = MEM[2208] + MEM[2286];
assign MEM[3810] = MEM[2209] + MEM[2227];
assign MEM[3811] = MEM[2209] + MEM[2248];
assign MEM[3812] = MEM[2210] + MEM[2333];
assign MEM[3813] = MEM[2216] + MEM[2298];
assign MEM[3814] = MEM[2219] + MEM[2235];
assign MEM[3815] = MEM[2221] + MEM[2238];
assign MEM[3816] = MEM[2222] + MEM[2232];
assign MEM[3817] = MEM[2222] + MEM[2236];
assign MEM[3818] = MEM[2225] + MEM[2254];
assign MEM[3819] = MEM[2227] + MEM[2394];
assign MEM[3820] = MEM[2230] + MEM[2276];
assign MEM[3821] = MEM[2231] + MEM[2321];
assign MEM[3822] = MEM[2232] + MEM[2254];
assign MEM[3823] = MEM[2235] + MEM[2274];
assign MEM[3824] = MEM[2236] + MEM[2311];
assign MEM[3825] = MEM[2237] + MEM[2286];
assign MEM[3826] = MEM[2238] + MEM[2278];
assign MEM[3827] = MEM[2239] + MEM[2340];
assign MEM[3828] = MEM[2240] + MEM[2241];
assign MEM[3829] = MEM[2241] + MEM[2304];
assign MEM[3830] = MEM[2243] + MEM[2267];
assign MEM[3831] = MEM[2244] + MEM[2292];
assign MEM[3832] = MEM[2244] + MEM[2332];
assign MEM[3833] = MEM[2245] + MEM[2258];
assign MEM[3834] = MEM[2245] + MEM[2321];
assign MEM[3835] = MEM[2247] + MEM[2306];
assign MEM[3836] = MEM[2248] + MEM[2301];
assign MEM[3837] = MEM[2252] + MEM[2281];
assign MEM[3838] = MEM[2252] + MEM[2284];
assign MEM[3839] = MEM[2256] + MEM[2258];
assign MEM[3840] = MEM[2256] + MEM[2320];
assign MEM[3841] = MEM[2257] + MEM[2273];
assign MEM[3842] = MEM[2257] + MEM[2359];
assign MEM[3843] = MEM[2262] + MEM[2275];
assign MEM[3844] = MEM[2266] + MEM[2291];
assign MEM[3845] = MEM[2266] + MEM[2402];
assign MEM[3846] = MEM[2270] + MEM[2272];
assign MEM[3847] = MEM[2270] + MEM[2309];
assign MEM[3848] = MEM[2271] + MEM[2330];
assign MEM[3849] = MEM[2271] + MEM[2342];
assign MEM[3850] = MEM[2272] + MEM[2450];
assign MEM[3851] = MEM[2273] + MEM[2301];
assign MEM[3852] = MEM[2274] + MEM[2349];
assign MEM[3853] = MEM[2276] + MEM[2281];
assign MEM[3854] = MEM[2277] + MEM[2279];
assign MEM[3855] = MEM[2277] + MEM[2280];
assign MEM[3856] = MEM[2278] + MEM[2307];
assign MEM[3857] = MEM[2279] + MEM[2437];
assign MEM[3858] = MEM[2280] + MEM[2285];
assign MEM[3859] = MEM[2283] + MEM[2304];
assign MEM[3860] = MEM[2290] + MEM[2331];
assign MEM[3861] = MEM[2290] + MEM[2372];
assign MEM[3862] = MEM[2291] + MEM[2370];
assign MEM[3863] = MEM[2293] + MEM[2308];
assign MEM[3864] = MEM[2293] + MEM[2363];
assign MEM[3865] = MEM[2297] + MEM[2369];
assign MEM[3866] = MEM[2298] + MEM[2306];
assign MEM[3867] = MEM[2307] + MEM[2422];
assign MEM[3868] = MEM[2308] + MEM[2344];
assign MEM[3869] = MEM[2309] + MEM[2327];
assign MEM[3870] = MEM[2310] + MEM[2327];
assign MEM[3871] = MEM[2311] + MEM[2356];
assign MEM[3872] = MEM[2313] + MEM[2328];
assign MEM[3873] = MEM[2313] + MEM[2335];
assign MEM[3874] = MEM[2314] + MEM[2331];
assign MEM[3875] = MEM[2314] + MEM[2349];
assign MEM[3876] = MEM[2315] + MEM[2323];
assign MEM[3877] = MEM[2315] + MEM[2517];
assign MEM[3878] = MEM[2317] + MEM[2319];
assign MEM[3879] = MEM[2317] + MEM[2332];
assign MEM[3880] = MEM[2318] + MEM[2361];
assign MEM[3881] = MEM[2318] + MEM[2420];
assign MEM[3882] = MEM[2319] + MEM[2389];
assign MEM[3883] = MEM[2320] + MEM[2358];
assign MEM[3884] = MEM[2323] + MEM[2388];
assign MEM[3885] = MEM[2325] + MEM[2339];
assign MEM[3886] = MEM[2325] + MEM[2465];
assign MEM[3887] = MEM[2328] + MEM[2362];
assign MEM[3888] = MEM[2330] + MEM[2410];
assign MEM[3889] = MEM[2333] + MEM[2525];
assign MEM[3890] = MEM[2335] + MEM[2348];
assign MEM[3891] = MEM[2336] + MEM[2375];
assign MEM[3892] = MEM[2336] + MEM[2413];
assign MEM[3893] = MEM[2339] + MEM[2391];
assign MEM[3894] = MEM[2340] + MEM[2447];
assign MEM[3895] = MEM[2341] + MEM[2351];
assign MEM[3896] = MEM[2341] + MEM[2354];
assign MEM[3897] = MEM[2342] + MEM[2377];
assign MEM[3898] = MEM[2343] + MEM[2388];
assign MEM[3899] = MEM[2344] + MEM[2354];
assign MEM[3900] = MEM[2347] + MEM[2350];
assign MEM[3901] = MEM[2348] + MEM[2395];
assign MEM[3902] = MEM[2350] + MEM[2351];
assign MEM[3903] = MEM[2355] + MEM[2424];
assign MEM[3904] = MEM[2355] + MEM[2491];
assign MEM[3905] = MEM[2356] + MEM[2436];
assign MEM[3906] = MEM[2357] + MEM[2362];
assign MEM[3907] = MEM[2357] + MEM[2448];
assign MEM[3908] = MEM[2358] + MEM[2375];
assign MEM[3909] = MEM[2359] + MEM[2387];
assign MEM[3910] = MEM[2360] + MEM[2366];
assign MEM[3911] = MEM[2361] + MEM[2569];
assign MEM[3912] = MEM[2363] + MEM[2371];
assign MEM[3913] = MEM[2366] + MEM[2455];
assign MEM[3914] = MEM[2369] + MEM[2444];
assign MEM[3915] = MEM[2370] + MEM[2389];
assign MEM[3916] = MEM[2371] + MEM[2374];
assign MEM[3917] = MEM[2372] + MEM[2380];
assign MEM[3918] = MEM[2374] + MEM[2403];
assign MEM[3919] = MEM[2377] + MEM[2393];
assign MEM[3920] = MEM[2378] + MEM[2382];
assign MEM[3921] = MEM[2378] + MEM[2449];
assign MEM[3922] = MEM[2379] + MEM[2405];
assign MEM[3923] = MEM[2379] + MEM[2500];
assign MEM[3924] = MEM[2380] + MEM[2495];
assign MEM[3925] = MEM[2382] + MEM[2479];
assign MEM[3926] = MEM[2384] + MEM[2391];
assign MEM[3927] = MEM[2384] + MEM[2614];
assign MEM[3928] = MEM[2386] + MEM[2413];
assign MEM[3929] = MEM[2386] + MEM[2414];
assign MEM[3930] = MEM[2387] + MEM[2405];
assign MEM[3931] = MEM[2392] + MEM[2393];
assign MEM[3932] = MEM[2392] + MEM[2471];
assign MEM[3933] = MEM[2394] + MEM[2429];
assign MEM[3934] = MEM[2395] + MEM[2421];
assign MEM[3935] = MEM[2402] + MEM[2414];
assign MEM[3936] = MEM[2403] + MEM[2468];
assign MEM[3937] = MEM[2407] + MEM[2432];
assign MEM[3938] = MEM[2407] + MEM[2497];
assign MEM[3939] = MEM[2410] + MEM[2492];
assign MEM[3940] = MEM[2412] + MEM[2420];
assign MEM[3941] = MEM[2412] + MEM[2461];
assign MEM[3942] = MEM[2419] + MEM[2475];
assign MEM[3943] = MEM[2421] + MEM[2434];
assign MEM[3944] = MEM[2422] + MEM[2554];
assign MEM[3945] = MEM[2424] + MEM[2430];
assign MEM[3946] = MEM[2429] + MEM[2455];
assign MEM[3947] = MEM[2430] + MEM[2438];
assign MEM[3948] = MEM[2431] + MEM[2437];
assign MEM[3949] = MEM[2431] + MEM[2440];
assign MEM[3950] = MEM[2432] + MEM[2444];
assign MEM[3951] = MEM[2433] + MEM[2500];
assign MEM[3952] = MEM[2433] + MEM[2566];
assign MEM[3953] = MEM[2434] + MEM[2521];
assign MEM[3954] = MEM[2436] + MEM[2482];
assign MEM[3955] = MEM[2438] + MEM[2471];
assign MEM[3956] = MEM[2439] + MEM[2489];
assign MEM[3957] = MEM[2439] + MEM[2512];
assign MEM[3958] = MEM[2440] + MEM[2449];
assign MEM[3959] = MEM[2441] + MEM[2459];
assign MEM[3960] = MEM[2441] + MEM[2587];
assign MEM[3961] = MEM[2443] + MEM[2483];
assign MEM[3962] = MEM[2443] + MEM[2511];
assign MEM[3963] = MEM[2447] + MEM[2457];
assign MEM[3964] = MEM[2448] + MEM[2467];
assign MEM[3965] = MEM[2450] + MEM[2488];
assign MEM[3966] = MEM[2451] + MEM[2463];
assign MEM[3967] = MEM[2451] + MEM[2511];
assign MEM[3968] = MEM[2456] + MEM[2469];
assign MEM[3969] = MEM[2456] + MEM[2476];
assign MEM[3970] = MEM[2457] + MEM[2463];
assign MEM[3971] = MEM[2459] + MEM[2566];
assign MEM[3972] = MEM[2461] + MEM[2468];
assign MEM[3973] = MEM[2464] + MEM[2491];
assign MEM[3974] = MEM[2464] + MEM[2504];
assign MEM[3975] = MEM[2465] + MEM[2543];
assign MEM[3976] = MEM[2467] + MEM[2497];
assign MEM[3977] = MEM[2469] + MEM[2472];
assign MEM[3978] = MEM[2470] + MEM[2485];
assign MEM[3979] = MEM[2470] + MEM[2493];
assign MEM[3980] = MEM[2472] + MEM[2485];
assign MEM[3981] = MEM[2475] + MEM[2498];
assign MEM[3982] = MEM[2476] + MEM[2532];
assign MEM[3983] = MEM[2478] + MEM[2514];
assign MEM[3984] = MEM[2478] + MEM[2540];
assign MEM[3985] = MEM[2479] + MEM[2498];
assign MEM[3986] = MEM[2482] + MEM[2539];
assign MEM[3987] = MEM[2483] + MEM[2510];
assign MEM[3988] = MEM[2484] + MEM[2541];
assign MEM[3989] = MEM[2484] + MEM[2565];
assign MEM[3990] = MEM[2487] + MEM[2519];
assign MEM[3991] = MEM[2487] + MEM[2537];
assign MEM[3992] = MEM[2488] + MEM[2593];
assign MEM[3993] = MEM[2489] + MEM[2493];
assign MEM[3994] = MEM[2492] + MEM[2522];
assign MEM[3995] = MEM[2495] + MEM[2551];
assign MEM[3996] = MEM[2496] + MEM[2533];
assign MEM[3997] = MEM[2496] + MEM[2567];
assign MEM[3998] = MEM[2504] + MEM[2536];
assign MEM[3999] = MEM[2507] + MEM[2541];
assign MEM[4000] = MEM[2507] + MEM[2701];
assign MEM[4001] = MEM[2508] + MEM[2512];
assign MEM[4002] = MEM[2508] + MEM[2518];
assign MEM[4003] = MEM[2509] + MEM[2533];
assign MEM[4004] = MEM[2509] + MEM[2549];
assign MEM[4005] = MEM[2510] + MEM[2625];
assign MEM[4006] = MEM[2514] + MEM[2550];
assign MEM[4007] = MEM[2515] + MEM[2555];
assign MEM[4008] = MEM[2515] + MEM[2570];
assign MEM[4009] = MEM[2517] + MEM[2546];
assign MEM[4010] = MEM[2518] + MEM[2583];
assign MEM[4011] = MEM[2519] + MEM[2571];
assign MEM[4012] = MEM[2521] + MEM[2585];
assign MEM[4013] = MEM[2522] + MEM[2534];
assign MEM[4014] = MEM[2523] + MEM[2529];
assign MEM[4015] = MEM[2523] + MEM[2589];
assign MEM[4016] = MEM[2525] + MEM[2593];
assign MEM[4017] = MEM[2529] + MEM[2573];
assign MEM[4018] = MEM[2532] + MEM[2556];
assign MEM[4019] = MEM[2534] + MEM[2549];
assign MEM[4020] = MEM[2536] + MEM[2557];
assign MEM[4021] = MEM[2537] + MEM[2616];
assign MEM[4022] = MEM[2539] + MEM[2575];
assign MEM[4023] = MEM[2540] + MEM[2576];
assign MEM[4024] = MEM[2542] + MEM[2545];
assign MEM[4025] = MEM[2542] + MEM[2625];
assign MEM[4026] = MEM[2543] + MEM[2560];
assign MEM[4027] = MEM[2545] + MEM[2551];
assign MEM[4028] = MEM[2546] + MEM[2618];
assign MEM[4029] = MEM[2548] + MEM[2588];
assign MEM[4030] = MEM[2548] + MEM[2612];
assign MEM[4031] = MEM[2550] + MEM[2579];
assign MEM[4032] = MEM[2553] + MEM[2555];
assign MEM[4033] = MEM[2553] + MEM[2602];
assign MEM[4034] = MEM[2554] + MEM[2656];
assign MEM[4035] = MEM[2556] + MEM[2564];
assign MEM[4036] = MEM[2557] + MEM[2574];
assign MEM[4037] = MEM[2560] + MEM[2567];
assign MEM[4038] = MEM[2561] + MEM[2617];
assign MEM[4039] = MEM[2561] + MEM[2650];
assign MEM[4040] = MEM[2562] + MEM[2595];
assign MEM[4041] = MEM[2562] + MEM[2644];
assign MEM[4042] = MEM[2564] + MEM[2599];
assign MEM[4043] = MEM[2565] + MEM[2685];
assign MEM[4044] = MEM[2569] + MEM[2684];
assign MEM[4045] = MEM[2570] + MEM[2573];
assign MEM[4046] = MEM[2571] + MEM[2579];
assign MEM[4047] = MEM[2574] + MEM[2651];
assign MEM[4048] = MEM[2575] + MEM[2601];
assign MEM[4049] = MEM[2576] + MEM[2594];
assign MEM[4050] = MEM[2580] + MEM[2583];
assign MEM[4051] = MEM[2580] + MEM[2610];
assign MEM[4052] = MEM[2582] + MEM[2586];
assign MEM[4053] = MEM[2582] + MEM[2607];
assign MEM[4054] = MEM[2584] + MEM[2634];
assign MEM[4055] = MEM[2584] + MEM[2636];
assign MEM[4056] = MEM[2585] + MEM[2652];
assign MEM[4057] = MEM[2586] + MEM[2592];
assign MEM[4058] = MEM[2587] + MEM[2710];
assign MEM[4059] = MEM[2588] + MEM[2683];
assign MEM[4060] = MEM[2589] + MEM[2591];
assign MEM[4061] = MEM[2590] + MEM[2748];
assign MEM[4062] = MEM[2590] + MEM[2751];
assign MEM[4063] = MEM[2591] + MEM[2697];
assign MEM[4064] = MEM[2592] + MEM[2598];
assign MEM[4065] = MEM[2594] + MEM[2680];
assign MEM[4066] = MEM[2595] + MEM[2635];
assign MEM[4067] = MEM[2596] + MEM[2642];
assign MEM[4068] = MEM[2596] + MEM[2669];
assign MEM[4069] = MEM[2598] + MEM[2613];
assign MEM[4070] = MEM[2599] + MEM[2733];
assign MEM[4071] = MEM[2601] + MEM[2617];
assign MEM[4072] = MEM[2602] + MEM[2669];
assign MEM[4073] = MEM[2603] + MEM[2638];
assign MEM[4074] = MEM[2603] + MEM[2699];
assign MEM[4075] = MEM[2606] + MEM[2612];
assign MEM[4076] = MEM[2606] + MEM[2645];
assign MEM[4077] = MEM[2607] + MEM[2699];
assign MEM[4078] = MEM[2610] + MEM[2754];
assign MEM[4079] = MEM[2613] + MEM[2619];
assign MEM[4080] = MEM[2614] + MEM[2616];
assign MEM[4081] = MEM[2618] + MEM[2751];
assign MEM[4082] = MEM[2619] + MEM[2678];
assign MEM[4083] = MEM[2624] + MEM[2631];
assign MEM[4084] = MEM[2624] + MEM[2639];
assign MEM[4085] = MEM[2626] + MEM[2651];
assign MEM[4086] = MEM[2626] + MEM[2678];
assign MEM[4087] = MEM[2628] + MEM[2645];
assign MEM[4088] = MEM[2628] + MEM[2763];
assign MEM[4089] = MEM[2631] + MEM[2674];
assign MEM[4090] = MEM[2632] + MEM[2640];
assign MEM[4091] = MEM[2632] + MEM[2750];
assign MEM[4092] = MEM[2633] + MEM[2664];
assign MEM[4093] = MEM[2633] + MEM[2680];
assign MEM[4094] = MEM[2634] + MEM[2642];
assign MEM[4095] = MEM[2635] + MEM[2638];
assign MEM[4096] = MEM[2636] + MEM[2664];
assign MEM[4097] = MEM[2639] + MEM[2679];
assign MEM[4098] = MEM[2640] + MEM[2701];
assign MEM[4099] = MEM[2644] + MEM[2708];
assign MEM[4100] = MEM[2649] + MEM[2685];
assign MEM[4101] = MEM[2649] + MEM[2687];
assign MEM[4102] = MEM[2650] + MEM[2656];
assign MEM[4103] = MEM[2652] + MEM[2688];
assign MEM[4104] = MEM[2653] + MEM[2691];
assign MEM[4105] = MEM[2653] + MEM[2697];
assign MEM[4106] = MEM[2654] + MEM[2670];
assign MEM[4107] = MEM[2654] + MEM[2735];
assign MEM[4108] = MEM[2658] + MEM[2684];
assign MEM[4109] = MEM[2658] + MEM[2715];
assign MEM[4110] = MEM[2659] + MEM[2663];
assign MEM[4111] = MEM[2659] + MEM[2711];
assign MEM[4112] = MEM[2663] + MEM[2740];
assign MEM[4113] = MEM[2665] + MEM[2666];
assign MEM[4114] = MEM[2665] + MEM[2719];
assign MEM[4115] = MEM[2666] + MEM[2714];
assign MEM[4116] = MEM[2668] + MEM[2720];
assign MEM[4117] = MEM[2668] + MEM[2775];
assign MEM[4118] = MEM[2670] + MEM[2681];
assign MEM[4119] = MEM[2674] + MEM[2677];
assign MEM[4120] = MEM[2677] + MEM[2733];
assign MEM[4121] = MEM[2679] + MEM[2762];
assign MEM[4122] = MEM[2681] + MEM[2718];
assign MEM[4123] = MEM[2682] + MEM[2707];
assign MEM[4124] = MEM[2682] + MEM[2708];
assign MEM[4125] = MEM[2683] + MEM[2780];
assign MEM[4126] = MEM[2687] + MEM[2702];
assign MEM[4127] = MEM[2688] + MEM[2690];
assign MEM[4128] = MEM[2690] + MEM[2722];
assign MEM[4129] = MEM[2691] + MEM[2702];
assign MEM[4130] = MEM[2692] + MEM[2741];
assign MEM[4131] = MEM[2692] + MEM[2759];
assign MEM[4132] = MEM[2693] + MEM[2725];
assign MEM[4133] = MEM[2693] + MEM[2737];
assign MEM[4134] = MEM[2704] + MEM[2724];
assign MEM[4135] = MEM[2704] + MEM[2744];
assign MEM[4136] = MEM[2707] + MEM[2760];
assign MEM[4137] = MEM[2709] + MEM[2710];
assign MEM[4138] = MEM[2709] + MEM[2725];
assign MEM[4139] = MEM[2711] + MEM[2746];
assign MEM[4140] = MEM[2714] + MEM[2732];
assign MEM[4141] = MEM[2715] + MEM[2717];
assign MEM[4142] = MEM[2716] + MEM[2736];
assign MEM[4143] = MEM[2716] + MEM[2759];
assign MEM[4144] = MEM[2717] + MEM[2723];
assign MEM[4145] = MEM[2718] + MEM[2743];
assign MEM[4146] = MEM[2719] + MEM[2737];
assign MEM[4147] = MEM[2720] + MEM[2731];
assign MEM[4148] = MEM[2722] + MEM[2750];
assign MEM[4149] = MEM[2723] + MEM[2742];
assign MEM[4150] = MEM[2724] + MEM[2758];
assign MEM[4151] = MEM[2727] + MEM[2735];
assign MEM[4152] = MEM[2727] + MEM[2801];
assign MEM[4153] = MEM[2728] + MEM[2776];
assign MEM[4154] = MEM[2728] + MEM[2813];
assign MEM[4155] = MEM[2731] + MEM[2739];
assign MEM[4156] = MEM[2732] + MEM[2743];
assign MEM[4157] = MEM[2734] + MEM[2784];
assign MEM[4158] = MEM[2734] + MEM[2794];
assign MEM[4159] = MEM[2736] + MEM[2796];
assign MEM[4160] = MEM[2738] + MEM[2749];
assign MEM[4161] = MEM[2738] + MEM[2791];
assign MEM[4162] = MEM[2739] + MEM[2754];
assign MEM[4163] = MEM[2740] + MEM[2809];
assign MEM[4164] = MEM[2741] + MEM[2773];
assign MEM[4165] = MEM[2742] + MEM[2803];
assign MEM[4166] = MEM[2744] + MEM[2777];
assign MEM[4167] = MEM[2745] + MEM[2746];
assign MEM[4168] = MEM[2745] + MEM[2793];
assign MEM[4169] = MEM[2747] + MEM[2752];
assign MEM[4170] = MEM[2747] + MEM[2793];
assign MEM[4171] = MEM[2748] + MEM[2796];
assign MEM[4172] = MEM[2749] + MEM[2776];
assign MEM[4173] = MEM[2752] + MEM[2797];
assign MEM[4174] = MEM[2753] + MEM[2806];
assign MEM[4175] = MEM[2753] + MEM[2809];
assign MEM[4176] = MEM[2755] + MEM[2756];
assign MEM[4177] = MEM[2755] + MEM[2780];
assign MEM[4178] = MEM[2756] + MEM[2823];
assign MEM[4179] = MEM[2757] + MEM[2763];
assign MEM[4180] = MEM[2757] + MEM[2806];
assign MEM[4181] = MEM[2758] + MEM[2781];
assign MEM[4182] = MEM[2760] + MEM[2835];
assign MEM[4183] = MEM[2761] + MEM[2767];
assign MEM[4184] = MEM[2761] + MEM[2773];
assign MEM[4185] = MEM[2762] + MEM[2772];
assign MEM[4186] = MEM[2764] + MEM[2767];
assign MEM[4187] = MEM[2764] + MEM[2857];
assign MEM[4188] = MEM[2765] + MEM[2772];
assign MEM[4189] = MEM[2765] + MEM[2778];
assign MEM[4190] = MEM[2766] + MEM[2781];
assign MEM[4191] = MEM[2766] + MEM[2879];
assign MEM[4192] = MEM[2768] + MEM[2787];
assign MEM[4193] = MEM[2768] + MEM[2807];
assign MEM[4194] = MEM[2770] + MEM[2779];
assign MEM[4195] = MEM[2770] + MEM[2811];
assign MEM[4196] = MEM[2771] + MEM[2778];
assign MEM[4197] = MEM[2771] + MEM[2782];
assign MEM[4198] = MEM[2774] + MEM[2783];
assign MEM[4199] = MEM[2774] + MEM[2856];
assign MEM[4200] = MEM[2775] + MEM[2918];
assign MEM[4201] = MEM[2777] + MEM[2820];
assign MEM[4202] = MEM[2779] + MEM[2785];
assign MEM[4203] = MEM[2782] + MEM[2787];
assign MEM[4204] = MEM[2783] + MEM[2808];
assign MEM[4205] = MEM[2784] + MEM[2816];
assign MEM[4206] = MEM[2785] + MEM[2805];
assign MEM[4207] = MEM[2786] + MEM[2802];
assign MEM[4208] = MEM[2786] + MEM[2823];
assign MEM[4209] = MEM[2788] + MEM[2804];
assign MEM[4210] = MEM[2788] + MEM[2824];
assign MEM[4211] = MEM[2789] + MEM[2800];
assign MEM[4212] = MEM[2789] + MEM[2942];
assign MEM[4213] = MEM[2790] + MEM[2804];
assign MEM[4214] = MEM[2790] + MEM[2869];
assign MEM[4215] = MEM[2791] + MEM[2814];
assign MEM[4216] = MEM[2792] + MEM[2795];
assign MEM[4217] = MEM[2792] + MEM[2885];
assign MEM[4218] = MEM[2794] + MEM[2812];
assign MEM[4219] = MEM[2795] + MEM[2801];
assign MEM[4220] = MEM[2797] + MEM[2848];
assign MEM[4221] = MEM[2798] + MEM[2812];
assign MEM[4222] = MEM[2798] + MEM[2836];
assign MEM[4223] = MEM[2799] + MEM[2817];
assign MEM[4224] = MEM[2799] + MEM[2831];
assign MEM[4225] = MEM[2800] + MEM[2825];
assign MEM[4226] = MEM[2802] + MEM[2830];
assign MEM[4227] = MEM[2803] + MEM[2815];
assign MEM[4228] = MEM[2805] + MEM[2842];
assign MEM[4229] = MEM[2807] + MEM[2833];
assign MEM[4230] = MEM[2808] + MEM[2911];
assign MEM[4231] = MEM[2810] + MEM[2816];
assign MEM[4232] = MEM[2810] + MEM[2832];
assign MEM[4233] = MEM[2811] + MEM[2820];
assign MEM[4234] = MEM[2813] + MEM[2876];
assign MEM[4235] = MEM[2814] + MEM[2831];
assign MEM[4236] = MEM[2815] + MEM[2873];
assign MEM[4237] = MEM[2817] + MEM[2844];
assign MEM[4238] = MEM[2818] + MEM[2822];
assign MEM[4239] = MEM[2818] + MEM[2825];
assign MEM[4240] = MEM[2821] + MEM[2840];
assign MEM[4241] = MEM[2821] + MEM[2859];
assign MEM[4242] = MEM[2822] + MEM[2830];
assign MEM[4243] = MEM[2824] + MEM[2835];
assign MEM[4244] = MEM[2826] + MEM[2845];
assign MEM[4245] = MEM[2826] + MEM[2891];
assign MEM[4246] = MEM[2827] + MEM[2849];
assign MEM[4247] = MEM[2827] + MEM[2851];
assign MEM[4248] = MEM[2828] + MEM[2846];
assign MEM[4249] = MEM[2828] + MEM[2858];
assign MEM[4250] = MEM[2829] + MEM[2839];
assign MEM[4251] = MEM[2829] + MEM[2866];
assign MEM[4252] = MEM[2832] + MEM[2864];
assign MEM[4253] = MEM[2833] + MEM[2834];
assign MEM[4254] = MEM[2834] + MEM[2847];
assign MEM[4255] = MEM[2836] + MEM[2865];
assign MEM[4256] = MEM[2837] + MEM[2838];
assign MEM[4257] = MEM[2837] + MEM[2884];
assign MEM[4258] = MEM[2838] + MEM[2888];
assign MEM[4259] = MEM[2839] + MEM[2841];
assign MEM[4260] = MEM[2840] + MEM[2884];
assign MEM[4261] = MEM[2841] + MEM[2862];
assign MEM[4262] = MEM[2842] + MEM[2937];
assign MEM[4263] = MEM[2843] + MEM[2860];
assign MEM[4264] = MEM[2843] + MEM[2881];
assign MEM[4265] = MEM[2844] + MEM[2846];
assign MEM[4266] = MEM[2845] + MEM[2899];
assign MEM[4267] = MEM[2847] + MEM[2985];
assign MEM[4268] = MEM[2848] + MEM[2945];
assign MEM[4269] = MEM[2849] + MEM[2883];
assign MEM[4270] = MEM[2850] + MEM[2876];
assign MEM[4271] = MEM[2850] + MEM[2922];
assign MEM[4272] = MEM[2851] + MEM[3004];
assign MEM[4273] = MEM[2852] + MEM[2853];
assign MEM[4274] = MEM[2852] + MEM[2861];
assign MEM[4275] = MEM[2853] + MEM[2871];
assign MEM[4276] = MEM[2854] + MEM[2862];
assign MEM[4277] = MEM[2854] + MEM[2917];
assign MEM[4278] = MEM[2855] + MEM[2877];
assign MEM[4279] = MEM[2855] + MEM[2907];
assign MEM[4280] = MEM[2856] + MEM[2898];
assign MEM[4281] = MEM[2857] + MEM[2887];
assign MEM[4282] = MEM[2858] + MEM[2870];
assign MEM[4283] = MEM[2859] + MEM[2990];
assign MEM[4284] = MEM[2860] + MEM[2963];
assign MEM[4285] = MEM[2861] + MEM[2927];
assign MEM[4286] = MEM[2863] + MEM[2940];
assign MEM[4287] = MEM[2863] + MEM[2949];
assign MEM[4288] = MEM[2864] + MEM[2872];
assign MEM[4289] = MEM[2865] + MEM[2915];
assign MEM[4290] = MEM[2866] + MEM[2931];
assign MEM[4291] = MEM[2867] + MEM[2871];
assign MEM[4292] = MEM[2867] + MEM[2881];
assign MEM[4293] = MEM[2868] + MEM[2872];
assign MEM[4294] = MEM[2868] + MEM[2916];
assign MEM[4295] = MEM[2869] + MEM[2939];
assign MEM[4296] = MEM[2870] + MEM[2971];
assign MEM[4297] = MEM[2873] + MEM[2894];
assign MEM[4298] = MEM[2874] + MEM[2878];
assign MEM[4299] = MEM[2874] + MEM[2936];
assign MEM[4300] = MEM[2875] + MEM[2895];
assign MEM[4301] = MEM[2875] + MEM[2956];
assign MEM[4302] = MEM[2877] + MEM[2886];
assign MEM[4303] = MEM[2878] + MEM[2919];
assign MEM[4304] = MEM[2879] + MEM[3174];
assign MEM[4305] = MEM[2880] + MEM[2929];
assign MEM[4306] = MEM[2880] + MEM[2953];
assign MEM[4307] = MEM[2882] + MEM[2890];
assign MEM[4308] = MEM[2882] + MEM[2896];
assign MEM[4309] = MEM[2883] + MEM[2959];
assign MEM[4310] = MEM[2885] + MEM[2944];
assign MEM[4311] = MEM[2886] + MEM[2938];
assign MEM[4312] = MEM[2889] + MEM[3011];
assign MEM[4313] = MEM[2892] + MEM[3057];
assign MEM[4314] = MEM[2893] + MEM[2948];
assign MEM[4315] = MEM[2897] + MEM[3101];
assign MEM[4316] = MEM[2900] + MEM[2957];
assign MEM[4317] = MEM[2901] + MEM[3005];
assign MEM[4318] = MEM[2902] + MEM[3026];
assign MEM[4319] = MEM[2903] + MEM[3031];
assign MEM[4320] = MEM[2904] + MEM[3039];
assign MEM[4321] = MEM[2905] + MEM[2969];
assign MEM[4322] = MEM[2906] + MEM[2999];
assign MEM[4323] = MEM[2908] + MEM[3038];
assign MEM[4324] = MEM[2909] + MEM[2954];
assign MEM[4325] = MEM[2910] + MEM[2992];
assign MEM[4326] = MEM[2912] + MEM[2983];
assign MEM[4327] = MEM[2913] + MEM[3046];
assign MEM[4328] = MEM[2914] + MEM[2997];
assign MEM[4329] = MEM[2920] + MEM[2930];
assign MEM[4330] = MEM[2921] + MEM[2962];
assign MEM[4331] = MEM[2923] + MEM[2950];
assign MEM[4332] = MEM[2924] + MEM[2935];
assign MEM[4333] = MEM[2925] + MEM[2984];
assign MEM[4334] = MEM[2926] + MEM[2974];
assign MEM[4335] = MEM[2928] + MEM[3047];
assign MEM[4336] = MEM[2932] + MEM[2966];
assign MEM[4337] = MEM[2933] + MEM[2961];
assign MEM[4338] = MEM[2934] + MEM[3003];
assign MEM[4339] = MEM[2941] + MEM[2987];
assign MEM[4340] = MEM[2943] + MEM[2981];
assign MEM[4341] = MEM[2946] + MEM[3032];
assign MEM[4342] = MEM[2947] + MEM[3118];
assign MEM[4343] = MEM[2951] + MEM[2986];
assign MEM[4344] = MEM[2952] + MEM[2989];
assign MEM[4345] = MEM[2955] + MEM[3014];
assign MEM[4346] = MEM[2958] + MEM[2988];
assign MEM[4347] = MEM[2960] + MEM[3007];
assign MEM[4348] = MEM[2964] + MEM[3052];
assign MEM[4349] = MEM[2965] + MEM[3110];
assign MEM[4350] = MEM[2967] + MEM[3009];
assign MEM[4351] = MEM[2968] + MEM[3055];
assign MEM[4352] = MEM[2970] + MEM[3017];
assign MEM[4353] = MEM[2972] + MEM[3024];
assign MEM[4354] = MEM[2973] + MEM[3021];
assign MEM[4355] = MEM[2975] + MEM[2982];
assign MEM[4356] = MEM[2976] + MEM[3030];
assign MEM[4357] = MEM[2977] + MEM[3015];
assign MEM[4358] = MEM[2978] + MEM[3054];
assign MEM[4359] = MEM[2979] + MEM[3071];
assign MEM[4360] = MEM[2980] + MEM[3070];
assign MEM[4361] = MEM[2991] + MEM[3034];
assign MEM[4362] = MEM[2993] + MEM[3002];
assign MEM[4363] = MEM[2994] + MEM[2995];
assign MEM[4364] = MEM[2996] + MEM[3245];
assign MEM[4365] = MEM[2998] + MEM[3018];
assign MEM[4366] = MEM[3000] + MEM[3069];
assign MEM[4367] = MEM[3001] + MEM[3027];
assign MEM[4368] = MEM[3006] + MEM[3122];
assign MEM[4369] = MEM[3008] + MEM[3133];
assign MEM[4370] = MEM[3010] + MEM[3041];
assign MEM[4371] = MEM[3012] + MEM[3090];
assign MEM[4372] = MEM[3013] + MEM[3072];
assign MEM[4373] = MEM[3016] + MEM[3053];
assign MEM[4374] = MEM[3019] + MEM[3093];
assign MEM[4375] = MEM[3020] + MEM[3104];
assign MEM[4376] = MEM[3022] + MEM[3105];
assign MEM[4377] = MEM[3023] + MEM[3119];
assign MEM[4378] = MEM[3025] + MEM[3162];
assign MEM[4379] = MEM[3028] + MEM[3060];
assign MEM[4380] = MEM[3029] + MEM[3043];
assign MEM[4381] = MEM[3033] + MEM[3078];
assign MEM[4382] = MEM[3035] + MEM[3091];
assign MEM[4383] = MEM[3036] + MEM[3111];
assign MEM[4384] = MEM[3037] + MEM[3040];
assign MEM[4385] = MEM[3042] + MEM[3114];
assign MEM[4386] = MEM[3044] + MEM[3061];
assign MEM[4387] = MEM[3045] + MEM[3066];
assign MEM[4388] = MEM[3048] + MEM[3199];
assign MEM[4389] = MEM[3049] + MEM[3109];
assign MEM[4390] = MEM[3050] + MEM[3176];
assign MEM[4391] = MEM[3051] + MEM[3186];
assign MEM[4392] = MEM[3056] + MEM[3079];
assign MEM[4393] = MEM[3058] + MEM[3124];
assign MEM[4394] = MEM[3059] + MEM[3121];
assign MEM[4395] = MEM[3062] + MEM[3168];
assign MEM[4396] = MEM[3063] + MEM[3081];
assign MEM[4397] = MEM[3064] + MEM[3087];
assign MEM[4398] = MEM[3065] + MEM[3113];
assign MEM[4399] = MEM[3067] + MEM[3085];
assign MEM[4400] = MEM[3068] + MEM[3089];
assign MEM[4401] = MEM[3073] + MEM[3147];
assign MEM[4402] = MEM[3074] + MEM[3116];
assign MEM[4403] = MEM[3075] + MEM[3259];
assign MEM[4404] = MEM[3076] + MEM[3137];
assign MEM[4405] = MEM[3077] + MEM[3117];
assign MEM[4406] = MEM[3080] + MEM[3139];
assign MEM[4407] = MEM[3082] + MEM[3276];
assign MEM[4408] = MEM[3083] + MEM[3185];
assign MEM[4409] = MEM[3084] + MEM[3144];
assign MEM[4410] = MEM[3086] + MEM[3149];
assign MEM[4411] = MEM[3088] + MEM[3177];
assign MEM[4412] = MEM[3092] + MEM[3107];
assign MEM[4413] = MEM[3094] + MEM[3163];
assign MEM[4414] = MEM[3095] + MEM[3181];
assign MEM[4415] = MEM[3096] + MEM[3112];
assign MEM[4416] = MEM[3097] + MEM[3134];
assign MEM[4417] = MEM[3098] + MEM[3115];
assign MEM[4418] = MEM[3099] + MEM[3428];
assign MEM[4419] = MEM[3100] + MEM[3130];
assign MEM[4420] = MEM[3102] + MEM[3142];
assign MEM[4421] = MEM[3103] + MEM[3165];
assign MEM[4422] = MEM[3106] + MEM[3178];
assign MEM[4423] = MEM[3108] + MEM[3209];
assign MEM[4424] = MEM[3120] + MEM[3152];
assign MEM[4425] = MEM[3123] + MEM[3160];
assign MEM[4426] = MEM[3125] + MEM[3205];
assign MEM[4427] = MEM[3126] + MEM[3217];
assign MEM[4428] = MEM[3127] + MEM[3151];
assign MEM[4429] = MEM[3128] + MEM[3164];
assign MEM[4430] = MEM[3129] + MEM[3157];
assign MEM[4431] = MEM[3131] + MEM[3288];
assign MEM[4432] = MEM[3132] + MEM[3155];
assign MEM[4433] = MEM[3135] + MEM[3169];
assign MEM[4434] = MEM[3136] + MEM[3224];
assign MEM[4435] = MEM[3138] + MEM[3241];
assign MEM[4436] = MEM[3140] + MEM[3183];
assign MEM[4437] = MEM[3141] + MEM[3289];
assign MEM[4438] = MEM[3143] + MEM[3179];
assign MEM[4439] = MEM[3145] + MEM[3171];
assign MEM[4440] = MEM[3146] + MEM[3211];
assign MEM[4441] = MEM[3148] + MEM[3197];
assign MEM[4442] = MEM[3150] + MEM[3194];
assign MEM[4443] = MEM[3153] + MEM[3240];
assign MEM[4444] = MEM[3154] + MEM[3238];
assign MEM[4445] = MEM[3156] + MEM[3187];
assign MEM[4446] = MEM[3158] + MEM[3254];
assign MEM[4447] = MEM[3159] + MEM[3215];
assign MEM[4448] = MEM[3161] + MEM[3268];
assign MEM[4449] = MEM[3166] + MEM[3258];
assign MEM[4450] = MEM[3167] + MEM[3216];
assign MEM[4451] = MEM[3170] + MEM[3300];
assign MEM[4452] = MEM[3172] + MEM[3203];
assign MEM[4453] = MEM[3173] + MEM[3255];
assign MEM[4454] = MEM[3175] + MEM[3202];
assign MEM[4455] = MEM[3180] + MEM[3235];
assign MEM[4456] = MEM[3182] + MEM[3272];
assign MEM[4457] = MEM[3184] + MEM[3232];
assign MEM[4458] = MEM[3188] + MEM[3298];
assign MEM[4459] = MEM[3189] + MEM[3244];
assign MEM[4460] = MEM[3190] + MEM[3234];
assign MEM[4461] = MEM[3191] + MEM[3242];
assign MEM[4462] = MEM[3192] + MEM[3247];
assign MEM[4463] = MEM[3193] + MEM[3207];
assign MEM[4464] = MEM[3195] + MEM[3219];
assign MEM[4465] = MEM[3196] + MEM[3319];
assign MEM[4466] = MEM[3198] + MEM[3229];
assign MEM[4467] = MEM[3200] + MEM[3256];
assign MEM[4468] = MEM[3201] + MEM[3344];
assign MEM[4469] = MEM[3204] + MEM[3233];
assign MEM[4470] = MEM[3206] + MEM[3271];
assign MEM[4471] = MEM[3208] + MEM[3239];
assign MEM[4472] = MEM[3210] + MEM[3267];
assign MEM[4473] = MEM[3212] + MEM[3269];
assign MEM[4474] = MEM[3213] + MEM[3304];
assign MEM[4475] = MEM[3214] + MEM[3370];
assign MEM[4476] = MEM[3218] + MEM[3225];
assign MEM[4477] = MEM[3220] + MEM[3237];
assign MEM[4478] = MEM[3221] + MEM[3281];
assign MEM[4479] = MEM[3222] + MEM[3236];
assign MEM[4480] = MEM[3223] + MEM[3310];
assign MEM[4481] = MEM[3226] + MEM[3470];
assign MEM[4482] = MEM[3227] + MEM[3264];
assign MEM[4483] = MEM[3228] + MEM[3263];
assign MEM[4484] = MEM[3230] + MEM[3329];
assign MEM[4485] = MEM[3231] + MEM[3305];
assign MEM[4486] = MEM[3243] + MEM[3309];
assign MEM[4487] = MEM[3246] + MEM[3279];
assign MEM[4488] = MEM[3248] + MEM[3261];
assign MEM[4489] = MEM[3249] + MEM[3295];
assign MEM[4490] = MEM[3250] + MEM[3374];
assign MEM[4491] = MEM[3251] + MEM[3301];
assign MEM[4492] = MEM[3252] + MEM[3342];
assign MEM[4493] = MEM[3253] + MEM[3318];
assign MEM[4494] = MEM[3257] + MEM[3278];
assign MEM[4495] = MEM[3260] + MEM[3262];
assign MEM[4496] = MEM[3265] + MEM[3345];
assign MEM[4497] = MEM[3266] + MEM[3395];
assign MEM[4498] = MEM[3270] + MEM[3283];
assign MEM[4499] = MEM[3273] + MEM[3315];
assign MEM[4500] = MEM[3274] + MEM[3320];
assign MEM[4501] = MEM[3275] + MEM[3338];
assign MEM[4502] = MEM[3277] + MEM[3293];
assign MEM[4503] = MEM[3280] + MEM[3384];
assign MEM[4504] = MEM[3282] + MEM[3316];
assign MEM[4505] = MEM[3284] + MEM[3379];
assign MEM[4506] = MEM[3285] + MEM[3323];
assign MEM[4507] = MEM[3286] + MEM[3314];
assign MEM[4508] = MEM[3287] + MEM[3381];
assign MEM[4509] = MEM[3290] + MEM[3363];
assign MEM[4510] = MEM[3291] + MEM[3386];
assign MEM[4511] = MEM[3292] + MEM[3339];
assign MEM[4512] = MEM[3294] + MEM[3404];
assign MEM[4513] = MEM[3296] + MEM[3340];
assign MEM[4514] = MEM[3297] + MEM[3324];
assign MEM[4515] = MEM[3299] + MEM[3341];
assign MEM[4516] = MEM[3302] + MEM[3365];
assign MEM[4517] = MEM[3303] + MEM[3372];
assign MEM[4518] = MEM[3306] + MEM[3393];
assign MEM[4519] = MEM[3307] + MEM[3353];
assign MEM[4520] = MEM[3308] + MEM[3334];
assign MEM[4521] = MEM[3311] + MEM[3336];
assign MEM[4522] = MEM[3312] + MEM[3333];
assign MEM[4523] = MEM[3313] + MEM[3397];
assign MEM[4524] = MEM[3317] + MEM[3354];
assign MEM[4525] = MEM[3321] + MEM[3411];
assign MEM[4526] = MEM[3322] + MEM[3408];
assign MEM[4527] = MEM[3325] + MEM[3366];
assign MEM[4528] = MEM[3326] + MEM[3414];
assign MEM[4529] = MEM[3327] + MEM[3383];
assign MEM[4530] = MEM[3328] + MEM[3361];
assign MEM[4531] = MEM[3330] + MEM[3377];
assign MEM[4532] = MEM[3331] + MEM[3419];
assign MEM[4533] = MEM[3332] + MEM[3390];
assign MEM[4534] = MEM[3335] + MEM[3448];
assign MEM[4535] = MEM[3337] + MEM[3475];
assign MEM[4536] = MEM[3343] + MEM[3410];
assign MEM[4537] = MEM[3346] + MEM[3422];
assign MEM[4538] = MEM[3347] + MEM[3369];
assign MEM[4539] = MEM[3348] + MEM[3382];
assign MEM[4540] = MEM[3349] + MEM[3423];
assign MEM[4541] = MEM[3350] + MEM[3398];
assign MEM[4542] = MEM[3351] + MEM[3405];
assign MEM[4543] = MEM[3352] + MEM[3378];
assign MEM[4544] = MEM[3355] + MEM[3455];
assign MEM[4545] = MEM[3356] + MEM[3389];
assign MEM[4546] = MEM[3357] + MEM[3436];
assign MEM[4547] = MEM[3358] + MEM[3406];
assign MEM[4548] = MEM[3359] + MEM[3418];
assign MEM[4549] = MEM[3360] + MEM[3429];
assign MEM[4550] = MEM[3362] + MEM[3385];
assign MEM[4551] = MEM[3364] + MEM[3416];
assign MEM[4552] = MEM[3367] + MEM[3391];
assign MEM[4553] = MEM[3368] + MEM[3407];
assign MEM[4554] = MEM[3371] + MEM[3430];
assign MEM[4555] = MEM[3373] + MEM[3457];
assign MEM[4556] = MEM[3375] + MEM[3464];
assign MEM[4557] = MEM[3376] + MEM[3554];
assign MEM[4558] = MEM[3380] + MEM[3424];
assign MEM[4559] = MEM[3387] + MEM[3486];
assign MEM[4560] = MEM[3388] + MEM[3412];
assign MEM[4561] = MEM[3392] + MEM[3447];
assign MEM[4562] = MEM[3394] + MEM[3468];
assign MEM[4563] = MEM[3396] + MEM[3485];
assign MEM[4564] = MEM[3399] + MEM[3454];
assign MEM[4565] = MEM[3400] + MEM[3420];
assign MEM[4566] = MEM[3401] + MEM[3467];
assign MEM[4567] = MEM[3402] + MEM[3462];
assign MEM[4568] = MEM[3403] + MEM[3444];
assign MEM[4569] = MEM[3409] + MEM[3489];
assign MEM[4570] = MEM[3413] + MEM[3518];
assign MEM[4571] = MEM[3415] + MEM[3588];
assign MEM[4572] = MEM[3417] + MEM[3510];
assign MEM[4573] = MEM[3421] + MEM[3491];
assign MEM[4574] = MEM[3425] + MEM[3503];
assign MEM[4575] = MEM[3426] + MEM[3469];
assign MEM[4576] = MEM[3427] + MEM[3471];
assign MEM[4577] = MEM[3431] + MEM[3541];
assign MEM[4578] = MEM[3432] + MEM[3465];
assign MEM[4579] = MEM[3433] + MEM[3459];
assign MEM[4580] = MEM[3434] + MEM[3458];
assign MEM[4581] = MEM[3435] + MEM[3476];
assign MEM[4582] = MEM[3437] + MEM[3497];
assign MEM[4583] = MEM[3438] + MEM[3584];
assign MEM[4584] = MEM[3439] + MEM[3446];
assign MEM[4585] = MEM[3440] + MEM[3498];
assign MEM[4586] = MEM[3441] + MEM[3500];
assign MEM[4587] = MEM[3442] + MEM[3449];
assign MEM[4588] = MEM[3443] + MEM[3521];
assign MEM[4589] = MEM[3445] + MEM[3482];
assign MEM[4590] = MEM[3450] + MEM[3477];
assign MEM[4591] = MEM[3451] + MEM[3513];
assign MEM[4592] = MEM[3452] + MEM[3511];
assign MEM[4593] = MEM[3453] + MEM[3478];
assign MEM[4594] = MEM[3456] + MEM[3529];
assign MEM[4595] = MEM[3460] + MEM[3526];
assign MEM[4596] = MEM[3461] + MEM[3642];
assign MEM[4597] = MEM[3463] + MEM[3496];
assign MEM[4598] = MEM[3466] + MEM[3539];
assign MEM[4599] = MEM[3472] + MEM[3532];
assign MEM[4600] = MEM[3473] + MEM[3553];
assign MEM[4601] = MEM[3474] + MEM[3638];
assign MEM[4602] = MEM[3479] + MEM[3537];
assign MEM[4603] = MEM[3480] + MEM[3587];
assign MEM[4604] = MEM[3481] + MEM[3528];
assign MEM[4605] = MEM[3483] + MEM[3502];
assign MEM[4606] = MEM[3484] + MEM[3558];
assign MEM[4607] = MEM[3487] + MEM[3555];
assign MEM[4608] = MEM[3488] + MEM[3585];
assign MEM[4609] = MEM[3490] + MEM[3544];
assign MEM[4610] = MEM[3492] + MEM[3495];
assign MEM[4611] = MEM[3493] + MEM[3561];
assign MEM[4612] = MEM[3494] + MEM[3501];
assign MEM[4613] = MEM[3499] + MEM[3508];
assign MEM[4614] = MEM[3504] + MEM[3575];
assign MEM[4615] = MEM[3505] + MEM[3551];
assign MEM[4616] = MEM[3506] + MEM[3591];
assign MEM[4617] = MEM[3507] + MEM[3548];
assign MEM[4618] = MEM[3509] + MEM[3547];
assign MEM[4619] = MEM[3512] + MEM[3579];
assign MEM[4620] = MEM[3514] + MEM[3538];
assign MEM[4621] = MEM[3515] + MEM[3612];
assign MEM[4622] = MEM[3516] + MEM[3534];
assign MEM[4623] = MEM[3517] + MEM[3581];
assign MEM[4624] = MEM[3519] + MEM[3545];
assign MEM[4625] = MEM[3520] + MEM[3572];
assign MEM[4626] = MEM[3522] + MEM[3556];
assign MEM[4627] = MEM[3523] + MEM[3562];
assign MEM[4628] = MEM[3524] + MEM[3629];
assign MEM[4629] = MEM[3525] + MEM[3598];
assign MEM[4630] = MEM[3527] + MEM[3613];
assign MEM[4631] = MEM[3530] + MEM[3606];
assign MEM[4632] = MEM[3531] + MEM[3576];
assign MEM[4633] = MEM[3533] + MEM[3624];
assign MEM[4634] = MEM[3535] + MEM[3649];
assign MEM[4635] = MEM[3536] + MEM[3696];
assign MEM[4636] = MEM[3540] + MEM[3567];
assign MEM[4637] = MEM[3542] + MEM[3608];
assign MEM[4638] = MEM[3543] + MEM[3633];
assign MEM[4639] = MEM[3546] + MEM[3574];
assign MEM[4640] = MEM[3549] + MEM[3623];
assign MEM[4641] = MEM[3550] + MEM[3621];
assign MEM[4642] = MEM[3552] + MEM[3568];
assign MEM[4643] = MEM[3557] + MEM[3569];
assign MEM[4644] = MEM[3559] + MEM[3565];
assign MEM[4645] = MEM[3560] + MEM[3596];
assign MEM[4646] = MEM[3563] + MEM[3685];
assign MEM[4647] = MEM[3564] + MEM[3609];
assign MEM[4648] = MEM[3566] + MEM[3819];
assign MEM[4649] = MEM[3570] + MEM[3618];
assign MEM[4650] = MEM[3571] + MEM[3657];
assign MEM[4651] = MEM[3573] + MEM[3600];
assign MEM[4652] = MEM[3577] + MEM[3676];
assign MEM[4653] = MEM[3578] + MEM[3586];
assign MEM[4654] = MEM[3580] + MEM[3615];
assign MEM[4655] = MEM[3582] + MEM[3603];
assign MEM[4656] = MEM[3583] + MEM[3658];
assign MEM[4657] = MEM[3589] + MEM[3605];
assign MEM[4658] = MEM[3590] + MEM[3660];
assign MEM[4659] = MEM[3592] + MEM[3648];
assign MEM[4660] = MEM[3593] + MEM[3782];
assign MEM[4661] = MEM[3594] + MEM[3715];
assign MEM[4662] = MEM[3595] + MEM[3708];
assign MEM[4663] = MEM[3597] + MEM[3644];
assign MEM[4664] = MEM[3599] + MEM[3710];
assign MEM[4665] = MEM[3601] + MEM[3674];
assign MEM[4666] = MEM[3602] + MEM[3650];
assign MEM[4667] = MEM[3604] + MEM[3688];
assign MEM[4668] = MEM[3607] + MEM[3634];
assign MEM[4669] = MEM[3610] + MEM[3637];
assign MEM[4670] = MEM[3611] + MEM[3697];
assign MEM[4671] = MEM[3614] + MEM[3640];
assign MEM[4672] = MEM[3616] + MEM[3625];
assign MEM[4673] = MEM[3617] + MEM[3639];
assign MEM[4674] = MEM[3619] + MEM[3761];
assign MEM[4675] = MEM[3620] + MEM[3635];
assign MEM[4676] = MEM[3622] + MEM[3680];
assign MEM[4677] = MEM[3626] + MEM[3667];
assign MEM[4678] = MEM[3627] + MEM[3668];
assign MEM[4679] = MEM[3628] + MEM[3751];
assign MEM[4680] = MEM[3630] + MEM[3821];
assign MEM[4681] = MEM[3631] + MEM[3641];
assign MEM[4682] = MEM[3632] + MEM[3707];
assign MEM[4683] = MEM[3636] + MEM[3730];
assign MEM[4684] = MEM[3643] + MEM[3767];
assign MEM[4685] = MEM[3645] + MEM[3722];
assign MEM[4686] = MEM[3646] + MEM[3690];
assign MEM[4687] = MEM[3647] + MEM[3682];
assign MEM[4688] = MEM[3651] + MEM[3747];
assign MEM[4689] = MEM[3652] + MEM[3744];
assign MEM[4690] = MEM[3653] + MEM[3739];
assign MEM[4691] = MEM[3654] + MEM[3663];
assign MEM[4692] = MEM[3655] + MEM[3681];
assign MEM[4693] = MEM[3656] + MEM[3694];
assign MEM[4694] = MEM[3659] + MEM[3671];
assign MEM[4695] = MEM[3661] + MEM[3714];
assign MEM[4696] = MEM[3662] + MEM[3840];
assign MEM[4697] = MEM[3664] + MEM[3699];
assign MEM[4698] = MEM[3665] + MEM[3695];
assign MEM[4699] = MEM[3666] + MEM[3770];
assign MEM[4700] = MEM[3669] + MEM[3709];
assign MEM[4701] = MEM[3670] + MEM[3678];
assign MEM[4702] = MEM[3672] + MEM[3718];
assign MEM[4703] = MEM[3673] + MEM[3733];
assign MEM[4704] = MEM[3675] + MEM[3754];
assign MEM[4705] = MEM[3677] + MEM[3771];
assign MEM[4706] = MEM[3679] + MEM[3746];
assign MEM[4707] = MEM[3683] + MEM[3720];
assign MEM[4708] = MEM[3684] + MEM[3801];
assign MEM[4709] = MEM[3686] + MEM[3740];
assign MEM[4710] = MEM[3687] + MEM[3768];
assign MEM[4711] = MEM[3689] + MEM[3842];
assign MEM[4712] = MEM[3691] + MEM[3864];
assign MEM[4713] = MEM[3692] + MEM[3738];
assign MEM[4714] = MEM[3693] + MEM[3781];
assign MEM[4715] = MEM[3698] + MEM[3712];
assign MEM[4716] = MEM[3700] + MEM[3734];
assign MEM[4717] = MEM[3701] + MEM[3723];
assign MEM[4718] = MEM[3702] + MEM[3780];
assign MEM[4719] = MEM[3703] + MEM[3798];
assign MEM[4720] = MEM[3704] + MEM[3745];
assign MEM[4721] = MEM[3705] + MEM[3721];
assign MEM[4722] = MEM[3706] + MEM[3732];
assign MEM[4723] = MEM[3711] + MEM[3717];
assign MEM[4724] = MEM[3713] + MEM[3743];
assign MEM[4725] = MEM[3716] + MEM[3809];
assign MEM[4726] = MEM[3719] + MEM[3796];
assign MEM[4727] = MEM[3724] + MEM[3736];
assign MEM[4728] = MEM[3725] + MEM[3753];
assign MEM[4729] = MEM[3726] + MEM[3776];
assign MEM[4730] = MEM[3727] + MEM[3784];
assign MEM[4731] = MEM[3728] + MEM[3766];
assign MEM[4732] = MEM[3729] + MEM[3769];
assign MEM[4733] = MEM[3731] + MEM[3762];
assign MEM[4734] = MEM[3735] + MEM[3788];
assign MEM[4735] = MEM[3737] + MEM[3752];
assign MEM[4736] = MEM[3741] + MEM[3831];
assign MEM[4737] = MEM[3742] + MEM[3812];
assign MEM[4738] = MEM[3748] + MEM[3797];
assign MEM[4739] = MEM[3749] + MEM[3837];
assign MEM[4740] = MEM[3750] + MEM[3810];
assign MEM[4741] = MEM[3755] + MEM[3824];
assign MEM[4742] = MEM[3756] + MEM[3814];
assign MEM[4743] = MEM[3757] + MEM[3789];
assign MEM[4744] = MEM[3758] + MEM[3785];
assign MEM[4745] = MEM[3759] + MEM[3787];
assign MEM[4746] = MEM[3760] + MEM[3792];
assign MEM[4747] = MEM[3763] + MEM[3851];
assign MEM[4748] = MEM[3764] + MEM[3856];
assign MEM[4749] = MEM[3765] + MEM[3841];
assign MEM[4750] = MEM[3772] + MEM[3857];
assign MEM[4751] = MEM[3773] + MEM[3846];
assign MEM[4752] = MEM[3774] + MEM[3813];
assign MEM[4753] = MEM[3775] + MEM[3826];
assign MEM[4754] = MEM[3777] + MEM[3938];
assign MEM[4755] = MEM[3778] + MEM[3873];
assign MEM[4756] = MEM[3779] + MEM[3811];
assign MEM[4757] = MEM[3783] + MEM[3817];
assign MEM[4758] = MEM[3786] + MEM[3818];
assign MEM[4759] = MEM[3790] + MEM[3872];
assign MEM[4760] = MEM[3791] + MEM[3808];
assign MEM[4761] = MEM[3793] + MEM[3986];
assign MEM[4762] = MEM[3794] + MEM[3888];
assign MEM[4763] = MEM[3795] + MEM[3900];
assign MEM[4764] = MEM[3799] + MEM[3852];
assign MEM[4765] = MEM[3800] + MEM[3984];
assign MEM[4766] = MEM[3802] + MEM[3959];
assign MEM[4767] = MEM[3803] + MEM[3843];
assign MEM[4768] = MEM[3804] + MEM[3839];
assign MEM[4769] = MEM[3805] + MEM[3862];
assign MEM[4770] = MEM[3806] + MEM[3901];
assign MEM[4771] = MEM[3807] + MEM[3827];
assign MEM[4772] = MEM[3815] + MEM[3956];
assign MEM[4773] = MEM[3816] + MEM[3874];
assign MEM[4774] = MEM[3820] + MEM[3883];
assign MEM[4775] = MEM[3822] + MEM[3855];
assign MEM[4776] = MEM[3823] + MEM[3853];
assign MEM[4777] = MEM[3825] + MEM[3903];
assign MEM[4778] = MEM[3828] + MEM[3866];
assign MEM[4779] = MEM[3829] + MEM[3892];
assign MEM[4780] = MEM[3830] + MEM[3847];
assign MEM[4781] = MEM[3832] + MEM[4008];
assign MEM[4782] = MEM[3833] + MEM[3879];
assign MEM[4783] = MEM[3834] + MEM[3918];
assign MEM[4784] = MEM[3835] + MEM[3876];
assign MEM[4785] = MEM[3836] + MEM[3935];
assign MEM[4786] = MEM[3838] + MEM[3878];
assign MEM[4787] = MEM[3844] + MEM[3867];
assign MEM[4788] = MEM[3845] + MEM[3988];
assign MEM[4789] = MEM[3848] + MEM[3895];
assign MEM[4790] = MEM[3849] + MEM[3925];
assign MEM[4791] = MEM[3850] + MEM[3982];
assign MEM[4792] = MEM[3854] + MEM[3877];
assign MEM[4793] = MEM[3858] + MEM[3896];
assign MEM[4794] = MEM[3859] + MEM[3947];
assign MEM[4795] = MEM[3860] + MEM[3893];
assign MEM[4796] = MEM[3861] + MEM[3952];
assign MEM[4797] = MEM[3863] + MEM[3904];
assign MEM[4798] = MEM[3865] + MEM[3915];
assign MEM[4799] = MEM[3868] + MEM[3945];
assign MEM[4800] = MEM[3869] + MEM[3941];
assign MEM[4801] = MEM[3870] + MEM[3908];
assign MEM[4802] = MEM[3871] + MEM[3994];
assign MEM[4803] = MEM[3875] + MEM[3920];
assign MEM[4804] = MEM[3880] + MEM[3921];
assign MEM[4805] = MEM[3881] + MEM[3964];
assign MEM[4806] = MEM[3882] + MEM[3976];
assign MEM[4807] = MEM[3884] + MEM[3960];
assign MEM[4808] = MEM[3885] + MEM[3924];
assign MEM[4809] = MEM[3886] + MEM[4005];
assign MEM[4810] = MEM[3887] + MEM[3979];
assign MEM[4811] = MEM[3889] + MEM[4030];
assign MEM[4812] = MEM[3890] + MEM[3905];
assign MEM[4813] = MEM[3891] + MEM[3927];
assign MEM[4814] = MEM[3894] + MEM[4011];
assign MEM[4815] = MEM[3897] + MEM[3990];
assign MEM[4816] = MEM[3898] + MEM[3932];
assign MEM[4817] = MEM[3899] + MEM[3911];
assign MEM[4818] = MEM[3902] + MEM[3928];
assign MEM[4819] = MEM[3906] + MEM[3957];
assign MEM[4820] = MEM[3907] + MEM[3966];
assign MEM[4821] = MEM[3909] + MEM[3974];
assign MEM[4822] = MEM[3910] + MEM[3950];
assign MEM[4823] = MEM[3912] + MEM[3981];
assign MEM[4824] = MEM[3913] + MEM[4003];
assign MEM[4825] = MEM[3914] + MEM[3972];
assign MEM[4826] = MEM[3916] + MEM[3919];
assign MEM[4827] = MEM[3917] + MEM[3973];
assign MEM[4828] = MEM[3922] + MEM[3968];
assign MEM[4829] = MEM[3923] + MEM[4053];
assign MEM[4830] = MEM[3926] + MEM[3987];
assign MEM[4831] = MEM[3929] + MEM[3942];
assign MEM[4832] = MEM[3930] + MEM[3944];
assign MEM[4833] = MEM[3931] + MEM[3937];
assign MEM[4834] = MEM[3933] + MEM[3954];
assign MEM[4835] = MEM[3934] + MEM[3955];
assign MEM[4836] = MEM[3936] + MEM[4004];
assign MEM[4837] = MEM[3939] + MEM[4015];
assign MEM[4838] = MEM[3940] + MEM[3951];
assign MEM[4839] = MEM[3943] + MEM[3970];
assign MEM[4840] = MEM[3946] + MEM[3980];
assign MEM[4841] = MEM[3948] + MEM[3971];
assign MEM[4842] = MEM[3949] + MEM[3965];
assign MEM[4843] = MEM[3953] + MEM[4105];
assign MEM[4844] = MEM[3958] + MEM[4020];
assign MEM[4845] = MEM[3961] + MEM[4027];
assign MEM[4846] = MEM[3962] + MEM[4043];
assign MEM[4847] = MEM[3963] + MEM[4028];
assign MEM[4848] = MEM[3967] + MEM[4021];
assign MEM[4849] = MEM[3969] + MEM[3991];
assign MEM[4850] = MEM[3975] + MEM[4050];
assign MEM[4851] = MEM[3977] + MEM[3993];
assign MEM[4852] = MEM[3978] + MEM[4056];
assign MEM[4853] = MEM[3983] + MEM[4038];
assign MEM[4854] = MEM[3985] + MEM[4017];
assign MEM[4855] = MEM[3989] + MEM[4118];
assign MEM[4856] = MEM[3992] + MEM[4111];
assign MEM[4857] = MEM[3995] + MEM[4033];
assign MEM[4858] = MEM[3996] + MEM[4061];
assign MEM[4859] = MEM[3997] + MEM[4048];
assign MEM[4860] = MEM[3998] + MEM[4075];
assign MEM[4861] = MEM[3999] + MEM[4103];
assign MEM[4862] = MEM[4000] + MEM[4145];
assign MEM[4863] = MEM[4001] + MEM[4068];
assign MEM[4864] = MEM[4002] + MEM[4013];
assign MEM[4865] = MEM[4006] + MEM[4051];
assign MEM[4866] = MEM[4007] + MEM[4067];
assign MEM[4867] = MEM[4009] + MEM[4101];
assign MEM[4868] = MEM[4010] + MEM[4079];
assign MEM[4869] = MEM[4012] + MEM[4084];
assign MEM[4870] = MEM[4014] + MEM[4040];
assign MEM[4871] = MEM[4016] + MEM[4096];
assign MEM[4872] = MEM[4018] + MEM[4091];
assign MEM[4873] = MEM[4019] + MEM[4057];
assign MEM[4874] = MEM[4022] + MEM[4055];
assign MEM[4875] = MEM[4023] + MEM[4097];
assign MEM[4876] = MEM[4024] + MEM[4074];
assign MEM[4877] = MEM[4025] + MEM[4088];
assign MEM[4878] = MEM[4026] + MEM[4093];
assign MEM[4879] = MEM[4029] + MEM[4107];
assign MEM[4880] = MEM[4031] + MEM[4083];
assign MEM[4881] = MEM[4032] + MEM[4036];
assign MEM[4882] = MEM[4034] + MEM[4119];
assign MEM[4883] = MEM[4035] + MEM[4071];
assign MEM[4884] = MEM[4037] + MEM[4052];
assign MEM[4885] = MEM[4039] + MEM[4142];
assign MEM[4886] = MEM[4041] + MEM[4100];
assign MEM[4887] = MEM[4042] + MEM[4077];
assign MEM[4888] = MEM[4044] + MEM[4134];
assign MEM[4889] = MEM[4045] + MEM[4117];
assign MEM[4890] = MEM[4046] + MEM[4072];
assign MEM[4891] = MEM[4047] + MEM[4115];
assign MEM[4892] = MEM[4049] + MEM[4086];
assign MEM[4893] = MEM[4054] + MEM[4156];
assign MEM[4894] = MEM[4058] + MEM[4216];
assign MEM[4895] = MEM[4059] + MEM[4168];
assign MEM[4896] = MEM[4060] + MEM[4102];
assign MEM[4897] = MEM[4062] + MEM[4177];
assign MEM[4898] = MEM[4063] + MEM[4136];
assign MEM[4899] = MEM[4064] + MEM[4104];
assign MEM[4900] = MEM[4065] + MEM[4132];
assign MEM[4901] = MEM[4066] + MEM[4306];
assign MEM[4902] = MEM[4069] + MEM[4188];
assign MEM[4903] = MEM[4070] + MEM[4158];
assign MEM[4904] = MEM[4073] + MEM[4129];
assign MEM[4905] = MEM[4076] + MEM[4112];
assign MEM[4906] = MEM[4078] + MEM[4181];
assign MEM[4907] = MEM[4080] + MEM[4089];
assign MEM[4908] = MEM[4081] + MEM[4195];
assign MEM[4909] = MEM[4082] + MEM[4141];
assign MEM[4910] = MEM[4085] + MEM[4116];
assign MEM[4911] = MEM[4087] + MEM[4106];
assign MEM[4912] = MEM[4090] + MEM[4114];
assign MEM[4913] = MEM[4092] + MEM[4138];
assign MEM[4914] = MEM[4094] + MEM[4164];
assign MEM[4915] = MEM[4095] + MEM[4125];
assign MEM[4916] = MEM[4098] + MEM[4201];
assign MEM[4917] = MEM[4099] + MEM[4171];
assign MEM[4918] = MEM[4108] + MEM[4133];
assign MEM[4919] = MEM[4109] + MEM[4163];
assign MEM[4920] = MEM[4110] + MEM[4131];
assign MEM[4921] = MEM[4113] + MEM[4124];
assign MEM[4922] = MEM[4120] + MEM[4199];
assign MEM[4923] = MEM[4121] + MEM[4303];
assign MEM[4924] = MEM[4122] + MEM[4162];
assign MEM[4925] = MEM[4123] + MEM[4214];
assign MEM[4926] = MEM[4126] + MEM[4144];
assign MEM[4927] = MEM[4127] + MEM[4192];
assign MEM[4928] = MEM[4128] + MEM[4178];
assign MEM[4929] = MEM[4130] + MEM[4173];
assign MEM[4930] = MEM[4135] + MEM[4167];
assign MEM[4931] = MEM[4137] + MEM[4146];
assign MEM[4932] = MEM[4139] + MEM[4187];
assign MEM[4933] = MEM[4140] + MEM[4204];
assign MEM[4934] = MEM[4143] + MEM[4243];
assign MEM[4935] = MEM[4147] + MEM[4159];
assign MEM[4936] = MEM[4148] + MEM[4186];
assign MEM[4937] = MEM[4149] + MEM[4218];
assign MEM[4938] = MEM[4150] + MEM[4230];
assign MEM[4939] = MEM[4151] + MEM[4175];
assign MEM[4940] = MEM[4152] + MEM[4238];
assign MEM[4941] = MEM[4153] + MEM[4210];
assign MEM[4942] = MEM[4154] + MEM[4235];
assign MEM[4943] = MEM[4155] + MEM[4212];
assign MEM[4944] = MEM[4157] + MEM[4245];
assign MEM[4945] = MEM[4160] + MEM[4211];
assign MEM[4946] = MEM[4161] + MEM[4249];
assign MEM[4947] = MEM[4165] + MEM[4237];
assign MEM[4948] = MEM[4166] + MEM[4240];
assign MEM[4949] = MEM[4169] + MEM[4221];
assign MEM[4950] = MEM[4170] + MEM[4219];
assign MEM[4951] = MEM[4172] + MEM[4255];
assign MEM[4952] = MEM[4174] + MEM[4233];
assign MEM[4953] = MEM[4176] + MEM[4256];
assign MEM[4954] = MEM[4179] + MEM[4209];
assign MEM[4955] = MEM[4180] + MEM[4232];
assign MEM[4956] = MEM[4182] + MEM[4281];
assign MEM[4957] = MEM[4183] + MEM[4231];
assign MEM[4958] = MEM[4184] + MEM[4206];
assign MEM[4959] = MEM[4185] + MEM[4285];
assign MEM[4960] = MEM[4189] + MEM[4261];
assign MEM[4961] = MEM[4190] + MEM[4225];
assign MEM[4962] = MEM[4191] + MEM[4324];
assign MEM[4963] = MEM[4193] + MEM[4236];
assign MEM[4964] = MEM[4194] + MEM[4203];
assign MEM[4965] = MEM[4196] + MEM[4229];
assign MEM[4966] = MEM[4197] + MEM[4208];
assign MEM[4967] = MEM[4198] + MEM[4226];
assign MEM[4968] = MEM[4200] + MEM[4364];
assign MEM[4969] = MEM[4202] + MEM[4258];
assign MEM[4970] = MEM[4205] + MEM[4260];
assign MEM[4971] = MEM[4207] + MEM[4283];
assign MEM[4972] = MEM[4213] + MEM[4251];
assign MEM[4973] = MEM[4215] + MEM[4239];
assign MEM[4974] = MEM[4217] + MEM[4319];
assign MEM[4975] = MEM[4220] + MEM[4323];
assign MEM[4976] = MEM[4222] + MEM[4268];
assign MEM[4977] = MEM[4223] + MEM[4309];
assign MEM[4978] = MEM[4224] + MEM[4278];
assign MEM[4979] = MEM[4227] + MEM[4242];
assign MEM[4980] = MEM[4228] + MEM[4299];
assign MEM[4981] = MEM[4234] + MEM[4305];
assign MEM[4982] = MEM[4241] + MEM[4292];
assign MEM[4983] = MEM[4244] + MEM[4284];
assign MEM[4984] = MEM[4246] + MEM[4279];
assign MEM[4985] = MEM[4247] + MEM[4290];
assign MEM[4986] = MEM[4248] + MEM[4328];
assign MEM[4987] = MEM[4250] + MEM[4264];
assign MEM[4988] = MEM[4252] + MEM[4339];
assign MEM[4989] = MEM[4253] + MEM[4257];
assign MEM[4990] = MEM[4254] + MEM[4302];
assign MEM[4991] = MEM[4259] + MEM[4274];
assign MEM[4992] = MEM[4262] + MEM[4359];
assign MEM[4993] = MEM[4263] + MEM[4289];
assign MEM[4994] = MEM[4265] + MEM[4275];
assign MEM[4995] = MEM[4266] + MEM[4336];
assign MEM[4996] = MEM[4267] + MEM[4400];
assign MEM[4997] = MEM[4269] + MEM[4314];
assign MEM[4998] = MEM[4270] + MEM[4335];
assign MEM[4999] = MEM[4271] + MEM[4371];
assign MEM[5000] = MEM[4272] + MEM[4382];
assign MEM[5001] = MEM[4273] + MEM[4315];
assign MEM[5002] = MEM[4276] + MEM[4391];
assign MEM[5003] = MEM[4277] + MEM[4372];
assign MEM[5004] = MEM[4280] + MEM[4358];
assign MEM[5005] = MEM[4282] + MEM[4307];
assign MEM[5006] = MEM[4286] + MEM[4342];
assign MEM[5007] = MEM[4287] + MEM[4361];
assign MEM[5008] = MEM[4288] + MEM[4377];
assign MEM[5009] = MEM[4291] + MEM[4340];
assign MEM[5010] = MEM[4293] + MEM[4313];
assign MEM[5011] = MEM[4294] + MEM[4379];
assign MEM[5012] = MEM[4295] + MEM[4375];
assign MEM[5013] = MEM[4296] + MEM[4421];
assign MEM[5014] = MEM[4297] + MEM[4341];
assign MEM[5015] = MEM[4298] + MEM[4304];
assign MEM[5016] = MEM[4300] + MEM[4356];
assign MEM[5017] = MEM[4301] + MEM[4357];
assign MEM[5018] = MEM[4308] + MEM[4329];
assign MEM[5019] = MEM[4310] + MEM[4351];
assign MEM[5020] = MEM[4311] + MEM[4344];
assign MEM[5021] = MEM[4312] + MEM[4390];
assign MEM[5022] = MEM[4316] + MEM[4368];
assign MEM[5023] = MEM[4317] + MEM[4388];
assign MEM[5024] = MEM[4318] + MEM[4420];
assign MEM[5025] = MEM[4320] + MEM[4412];
assign MEM[5026] = MEM[4321] + MEM[4387];
assign MEM[5027] = MEM[4322] + MEM[4393];
assign MEM[5028] = MEM[4325] + MEM[4398];
assign MEM[5029] = MEM[4326] + MEM[4386];
assign MEM[5030] = MEM[4327] + MEM[4402];
assign MEM[5031] = MEM[4330] + MEM[4354];
assign MEM[5032] = MEM[4331] + MEM[4417];
assign MEM[5033] = MEM[4332] + MEM[4363];
assign MEM[5034] = MEM[4333] + MEM[4380];
assign MEM[5035] = MEM[4334] + MEM[4366];
assign MEM[5036] = MEM[4337] + MEM[4370];
assign MEM[5037] = MEM[4338] + MEM[4407];
assign MEM[5038] = MEM[4343] + MEM[4397];
assign MEM[5039] = MEM[4345] + MEM[4477];
assign MEM[5040] = MEM[4346] + MEM[4381];
assign MEM[5041] = MEM[4347] + MEM[4374];
assign MEM[5042] = MEM[4348] + MEM[4396];
assign MEM[5043] = MEM[4349] + MEM[4449];
assign MEM[5044] = MEM[4350] + MEM[4411];
assign MEM[5045] = MEM[4352] + MEM[4432];
assign MEM[5046] = MEM[4353] + MEM[4414];
assign MEM[5047] = MEM[4355] + MEM[4369];
assign MEM[5048] = MEM[4360] + MEM[4405];
assign MEM[5049] = MEM[4362] + MEM[4383];
assign MEM[5050] = MEM[4365] + MEM[4406];
assign MEM[5051] = MEM[4367] + MEM[4430];
assign MEM[5052] = MEM[4373] + MEM[4404];
assign MEM[5053] = MEM[4376] + MEM[4443];
assign MEM[5054] = MEM[4378] + MEM[4510];
assign MEM[5055] = MEM[4384] + MEM[4416];
assign MEM[5056] = MEM[4385] + MEM[4440];
assign MEM[5057] = MEM[4389] + MEM[4446];
assign MEM[5058] = MEM[4392] + MEM[4429];
assign MEM[5059] = MEM[4394] + MEM[4452];
assign MEM[5060] = MEM[4395] + MEM[4456];
assign MEM[5061] = MEM[4399] + MEM[4435];
assign MEM[5062] = MEM[4401] + MEM[4460];
assign MEM[5063] = MEM[4403] + MEM[4528];
assign MEM[5064] = MEM[4408] + MEM[4494];
assign MEM[5065] = MEM[4409] + MEM[4457];
assign MEM[5066] = MEM[4410] + MEM[4462];
assign MEM[5067] = MEM[4413] + MEM[4472];
assign MEM[5068] = MEM[4415] + MEM[4493];
assign MEM[5069] = MEM[4418] + MEM[4594];
assign MEM[5070] = MEM[4419] + MEM[4444];
assign MEM[5071] = MEM[4422] + MEM[4484];
assign MEM[5072] = MEM[4423] + MEM[4517];
assign MEM[5073] = MEM[4424] + MEM[4448];
assign MEM[5074] = MEM[4425] + MEM[4461];
assign MEM[5075] = MEM[4426] + MEM[4489];
assign MEM[5076] = MEM[4427] + MEM[4487];
assign MEM[5077] = MEM[4428] + MEM[4470];
assign MEM[5078] = MEM[4431] + MEM[4520];
assign MEM[5079] = MEM[4433] + MEM[4469];
assign MEM[5080] = MEM[4434] + MEM[4509];
assign MEM[5081] = MEM[4436] + MEM[4485];
assign MEM[5082] = MEM[4437] + MEM[4560];
assign MEM[5083] = MEM[4438] + MEM[4466];
assign MEM[5084] = MEM[4439] + MEM[4500];
assign MEM[5085] = MEM[4441] + MEM[4488];
assign MEM[5086] = MEM[4442] + MEM[4495];
assign MEM[5087] = MEM[4445] + MEM[4526];
assign MEM[5088] = MEM[4447] + MEM[4503];
assign MEM[5089] = MEM[4450] + MEM[4478];
assign MEM[5090] = MEM[4451] + MEM[4548];
assign MEM[5091] = MEM[4453] + MEM[4525];
assign MEM[5092] = MEM[4454] + MEM[4475];
assign MEM[5093] = MEM[4455] + MEM[4508];
assign MEM[5094] = MEM[4458] + MEM[4539];
assign MEM[5095] = MEM[4459] + MEM[4521];
assign MEM[5096] = MEM[4463] + MEM[4505];
assign MEM[5097] = MEM[4464] + MEM[4491];
assign MEM[5098] = MEM[4465] + MEM[4587];
assign MEM[5099] = MEM[4467] + MEM[4515];
assign MEM[5100] = MEM[4468] + MEM[4595];
assign MEM[5101] = MEM[4471] + MEM[4498];
assign MEM[5102] = MEM[4473] + MEM[4513];
assign MEM[5103] = MEM[4474] + MEM[4568];
assign MEM[5104] = MEM[4476] + MEM[4518];
assign MEM[5105] = MEM[4479] + MEM[4490];
assign MEM[5106] = MEM[4480] + MEM[4544];
assign MEM[5107] = MEM[4481] + MEM[4638];
assign MEM[5108] = MEM[4482] + MEM[4504];
assign MEM[5109] = MEM[4483] + MEM[4564];
assign MEM[5110] = MEM[4486] + MEM[4529];
assign MEM[5111] = MEM[4492] + MEM[4627];
assign MEM[5112] = MEM[4496] + MEM[4566];
assign MEM[5113] = MEM[4497] + MEM[4572];
assign MEM[5114] = MEM[4499] + MEM[4538];
assign MEM[5115] = MEM[4501] + MEM[4567];
assign MEM[5116] = MEM[4502] + MEM[4562];
assign MEM[5117] = MEM[4506] + MEM[4558];
assign MEM[5118] = MEM[4507] + MEM[4543];
assign MEM[5119] = MEM[4511] + MEM[4550];
assign MEM[5120] = MEM[4512] + MEM[4584];
assign MEM[5121] = MEM[4514] + MEM[4537];
assign MEM[5122] = MEM[4516] + MEM[4608];
assign MEM[5123] = MEM[4519] + MEM[4578];
assign MEM[5124] = MEM[4522] + MEM[4547];
assign MEM[5125] = MEM[4523] + MEM[4580];
assign MEM[5126] = MEM[4524] + MEM[4641];
assign MEM[5127] = MEM[4527] + MEM[4585];
assign MEM[5128] = MEM[4530] + MEM[4569];
assign MEM[5129] = MEM[4531] + MEM[4577];
assign MEM[5130] = MEM[4532] + MEM[4579];
assign MEM[5131] = MEM[4533] + MEM[4576];
assign MEM[5132] = MEM[4534] + MEM[4614];
assign MEM[5133] = MEM[4535] + MEM[4708];
assign MEM[5134] = MEM[4536] + MEM[4581];
assign MEM[5135] = MEM[4540] + MEM[4605];
assign MEM[5136] = MEM[4541] + MEM[4570];
assign MEM[5137] = MEM[4542] + MEM[4583];
assign MEM[5138] = MEM[4545] + MEM[4632];
assign MEM[5139] = MEM[4546] + MEM[4625];
assign MEM[5140] = MEM[4549] + MEM[4612];
assign MEM[5141] = MEM[4551] + MEM[4599];
assign MEM[5142] = MEM[4552] + MEM[4573];
assign MEM[5143] = MEM[4553] + MEM[4596];
assign MEM[5144] = MEM[4554] + MEM[4657];
assign MEM[5145] = MEM[4555] + MEM[4607];
assign MEM[5146] = MEM[4556] + MEM[4618];
assign MEM[5147] = MEM[4557] + MEM[4645];
assign MEM[5148] = MEM[4559] + MEM[4628];
assign MEM[5149] = MEM[4561] + MEM[4609];
assign MEM[5150] = MEM[4563] + MEM[4620];
assign MEM[5151] = MEM[4565] + MEM[4610];
assign MEM[5152] = MEM[4571] + MEM[4670];
assign MEM[5153] = MEM[4574] + MEM[4658];
assign MEM[5154] = MEM[4575] + MEM[4611];
assign MEM[5155] = MEM[4582] + MEM[4622];
assign MEM[5156] = MEM[4586] + MEM[4644];
assign MEM[5157] = MEM[4588] + MEM[4643];
assign MEM[5158] = MEM[4589] + MEM[4660];
assign MEM[5159] = MEM[4590] + MEM[4676];
assign MEM[5160] = MEM[4591] + MEM[4636];
assign MEM[5161] = MEM[4592] + MEM[4652];
assign MEM[5162] = MEM[4593] + MEM[4655];
assign MEM[5163] = MEM[4597] + MEM[4629];
assign MEM[5164] = MEM[4598] + MEM[4671];
assign MEM[5165] = MEM[4600] + MEM[4675];
assign MEM[5166] = MEM[4601] + MEM[4704];
assign MEM[5167] = MEM[4602] + MEM[4648];
assign MEM[5168] = MEM[4603] + MEM[4724];
assign MEM[5169] = MEM[4604] + MEM[4650];
assign MEM[5170] = MEM[4606] + MEM[4685];
assign MEM[5171] = MEM[4613] + MEM[4642];
assign MEM[5172] = MEM[4615] + MEM[4656];
assign MEM[5173] = MEM[4616] + MEM[4692];
assign MEM[5174] = MEM[4617] + MEM[4693];
assign MEM[5175] = MEM[4619] + MEM[4705];
assign MEM[5176] = MEM[4621] + MEM[4706];
assign MEM[5177] = MEM[4623] + MEM[4662];
assign MEM[5178] = MEM[4624] + MEM[4672];
assign MEM[5179] = MEM[4626] + MEM[4683];
assign MEM[5180] = MEM[4630] + MEM[4694];
assign MEM[5181] = MEM[4631] + MEM[4679];
assign MEM[5182] = MEM[4633] + MEM[4734];
assign MEM[5183] = MEM[4634] + MEM[4699];
assign MEM[5184] = MEM[4635] + MEM[4751];
assign MEM[5185] = MEM[4637] + MEM[4747];
assign MEM[5186] = MEM[4639] + MEM[4661];
assign MEM[5187] = MEM[4640] + MEM[4723];
assign MEM[5188] = MEM[4646] + MEM[4721];
assign MEM[5189] = MEM[4647] + MEM[4702];
assign MEM[5190] = MEM[4649] + MEM[4727];
assign MEM[5191] = MEM[4651] + MEM[4725];
assign MEM[5192] = MEM[4653] + MEM[4689];
assign MEM[5193] = MEM[4654] + MEM[4680];
assign MEM[5194] = MEM[4659] + MEM[4755];
assign MEM[5195] = MEM[4663] + MEM[4712];
assign MEM[5196] = MEM[4664] + MEM[4735];
assign MEM[5197] = MEM[4665] + MEM[4741];
assign MEM[5198] = MEM[4666] + MEM[4740];
assign MEM[5199] = MEM[4667] + MEM[4713];
assign MEM[5200] = MEM[4668] + MEM[4739];
assign MEM[5201] = MEM[4669] + MEM[4749];
assign MEM[5202] = MEM[4673] + MEM[4710];
assign MEM[5203] = MEM[4674] + MEM[4785];
assign MEM[5204] = MEM[4677] + MEM[4711];
assign MEM[5205] = MEM[4678] + MEM[4722];
assign MEM[5206] = MEM[4681] + MEM[4716];
assign MEM[5207] = MEM[4682] + MEM[4744];
assign MEM[5208] = MEM[4684] + MEM[4776];
assign MEM[5209] = MEM[4686] + MEM[4754];
assign MEM[5210] = MEM[4687] + MEM[4731];
assign MEM[5211] = MEM[4688] + MEM[4750];
assign MEM[5212] = MEM[4690] + MEM[4758];
assign MEM[5213] = MEM[4691] + MEM[4718];
assign MEM[5214] = MEM[4695] + MEM[4763];
assign MEM[5215] = MEM[4696] + MEM[4807];
assign MEM[5216] = MEM[4697] + MEM[4729];
assign MEM[5217] = MEM[4698] + MEM[4760];
assign MEM[5218] = MEM[4700] + MEM[4730];
assign MEM[5219] = MEM[4701] + MEM[4714];
assign MEM[5220] = MEM[4703] + MEM[4775];
assign MEM[5221] = MEM[4707] + MEM[4752];
assign MEM[5222] = MEM[4709] + MEM[4771];
assign MEM[5223] = MEM[4715] + MEM[4732];
assign MEM[5224] = MEM[4717] + MEM[4737];
assign MEM[5225] = MEM[4719] + MEM[4800];
assign MEM[5226] = MEM[4720] + MEM[4757];
assign MEM[5227] = MEM[4726] + MEM[4779];
assign MEM[5228] = MEM[4728] + MEM[4778];
assign MEM[5229] = MEM[4733] + MEM[4777];
assign MEM[5230] = MEM[4736] + MEM[4805];
assign MEM[5231] = MEM[4738] + MEM[4787];
assign MEM[5232] = MEM[4742] + MEM[4780];
assign MEM[5233] = MEM[4743] + MEM[4822];
assign MEM[5234] = MEM[4745] + MEM[4806];
assign MEM[5235] = MEM[4746] + MEM[4783];
assign MEM[5236] = MEM[4748] + MEM[4803];
assign MEM[5237] = MEM[4753] + MEM[4795];
assign MEM[5238] = MEM[4756] + MEM[4794];
assign MEM[5239] = MEM[4759] + MEM[4813];
assign MEM[5240] = MEM[4761] + MEM[4883];
assign MEM[5241] = MEM[4762] + MEM[4847];
assign MEM[5242] = MEM[4764] + MEM[4818];
assign MEM[5243] = MEM[4765] + MEM[4904];
assign MEM[5244] = MEM[4766] + MEM[4860];
assign MEM[5245] = MEM[4767] + MEM[4819];
assign MEM[5246] = MEM[4768] + MEM[4804];
assign MEM[5247] = MEM[4769] + MEM[4834];
assign MEM[5248] = MEM[4770] + MEM[4864];
assign MEM[5249] = MEM[4772] + MEM[4858];
assign MEM[5250] = MEM[4773] + MEM[4811];
assign MEM[5251] = MEM[4774] + MEM[4823];
assign MEM[5252] = MEM[4781] + MEM[4903];
assign MEM[5253] = MEM[4782] + MEM[4814];
assign MEM[5254] = MEM[4784] + MEM[4815];
assign MEM[5255] = MEM[4786] + MEM[4817];
assign MEM[5256] = MEM[4788] + MEM[4900];
assign MEM[5257] = MEM[4789] + MEM[4825];
assign MEM[5258] = MEM[4790] + MEM[4869];
assign MEM[5259] = MEM[4791] + MEM[4884];
assign MEM[5260] = MEM[4792] + MEM[4872];
assign MEM[5261] = MEM[4793] + MEM[4867];
assign MEM[5262] = MEM[4796] + MEM[4896];
assign MEM[5263] = MEM[4797] + MEM[4859];
assign MEM[5264] = MEM[4798] + MEM[4833];
assign MEM[5265] = MEM[4799] + MEM[4932];
assign MEM[5266] = MEM[4801] + MEM[4851];
assign MEM[5267] = MEM[4802] + MEM[4891];
assign MEM[5268] = MEM[4808] + MEM[4874];
assign MEM[5269] = MEM[4809] + MEM[4910];
assign MEM[5270] = MEM[4810] + MEM[4865];
assign MEM[5271] = MEM[4812] + MEM[4844];
assign MEM[5272] = MEM[4816] + MEM[4856];
assign MEM[5273] = MEM[4820] + MEM[4886];
assign MEM[5274] = MEM[4821] + MEM[4861];
assign MEM[5275] = MEM[4824] + MEM[4882];
assign MEM[5276] = MEM[4826] + MEM[4837];
assign MEM[5277] = MEM[4827] + MEM[4868];
assign MEM[5278] = MEM[4828] + MEM[4855];
assign MEM[5279] = MEM[4829] + MEM[4907];
assign MEM[5280] = MEM[4830] + MEM[4890];
assign MEM[5281] = MEM[4831] + MEM[4928];
assign MEM[5282] = MEM[4832] + MEM[4887];
assign MEM[5283] = MEM[4835] + MEM[4853];
assign MEM[5284] = MEM[4836] + MEM[4885];
assign MEM[5285] = MEM[4838] + MEM[4876];
assign MEM[5286] = MEM[4839] + MEM[4850];
assign MEM[5287] = MEM[4840] + MEM[4857];
assign MEM[5288] = MEM[4841] + MEM[4909];
assign MEM[5289] = MEM[4842] + MEM[4879];
assign MEM[5290] = MEM[4843] + MEM[4937];
assign MEM[5291] = MEM[4845] + MEM[4893];
assign MEM[5292] = MEM[4846] + MEM[4953];
assign MEM[5293] = MEM[4848] + MEM[4916];
assign MEM[5294] = MEM[4849] + MEM[4898];
assign MEM[5295] = MEM[4852] + MEM[4940];
assign MEM[5296] = MEM[4854] + MEM[4899];
assign MEM[5297] = MEM[4862] + MEM[4977];
assign MEM[5298] = MEM[4863] + MEM[4930];
assign MEM[5299] = MEM[4866] + MEM[4951];
assign MEM[5300] = MEM[4870] + MEM[4906];
assign MEM[5301] = MEM[4871] + MEM[4922];
assign MEM[5302] = MEM[4873] + MEM[4919];
assign MEM[5303] = MEM[4875] + MEM[4935];
assign MEM[5304] = MEM[4877] + MEM[4966];
assign MEM[5305] = MEM[4878] + MEM[4976];
assign MEM[5306] = MEM[4880] + MEM[4924];
assign MEM[5307] = MEM[4881] + MEM[4895];
assign MEM[5308] = MEM[4888] + MEM[4946];
assign MEM[5309] = MEM[4889] + MEM[4978];
assign MEM[5310] = MEM[4892] + MEM[4925];
assign MEM[5311] = MEM[4894] + MEM[4975];
assign MEM[5312] = MEM[4897] + MEM[4988];
assign MEM[5313] = MEM[4901] + MEM[5042];
assign MEM[5314] = MEM[4902] + MEM[4979];
assign MEM[5315] = MEM[4905] + MEM[5025];
assign MEM[5316] = MEM[4908] + MEM[4989];
assign MEM[5317] = MEM[4911] + MEM[4931];
assign MEM[5318] = MEM[4912] + MEM[4950];
assign MEM[5319] = MEM[4913] + MEM[4962];
assign MEM[5320] = MEM[4914] + MEM[4968];
assign MEM[5321] = MEM[4915] + MEM[4971];
assign MEM[5322] = MEM[4917] + MEM[5020];
assign MEM[5323] = MEM[4918] + MEM[4963];
assign MEM[5324] = MEM[4920] + MEM[4964];
assign MEM[5325] = MEM[4921] + MEM[4943];
assign MEM[5326] = MEM[4923] + MEM[5043];
assign MEM[5327] = MEM[4926] + MEM[4944];
assign MEM[5328] = MEM[4927] + MEM[4980];
assign MEM[5329] = MEM[4929] + MEM[4982];
assign MEM[5330] = MEM[4933] + MEM[4990];
assign MEM[5331] = MEM[4934] + MEM[4992];
assign MEM[5332] = MEM[4936] + MEM[4972];
assign MEM[5333] = MEM[4938] + MEM[5047];
assign MEM[5334] = MEM[4939] + MEM[5001];
assign MEM[5335] = MEM[4941] + MEM[4995];
assign MEM[5336] = MEM[4942] + MEM[4993];
assign MEM[5337] = MEM[4945] + MEM[4997];
assign MEM[5338] = MEM[4947] + MEM[5004];
assign MEM[5339] = MEM[4948] + MEM[4996];
assign MEM[5340] = MEM[4949] + MEM[5024];
assign MEM[5341] = MEM[4952] + MEM[5035];
assign MEM[5342] = MEM[4954] + MEM[4994];
assign MEM[5343] = MEM[4955] + MEM[5027];
assign MEM[5344] = MEM[4956] + MEM[5034];
assign MEM[5345] = MEM[4957] + MEM[5012];
assign MEM[5346] = MEM[4958] + MEM[5010];
assign MEM[5347] = MEM[4959] + MEM[5040];
assign MEM[5348] = MEM[4960] + MEM[5011];
assign MEM[5349] = MEM[4961] + MEM[5007];
assign MEM[5350] = MEM[4965] + MEM[5013];
assign MEM[5351] = MEM[4967] + MEM[5000];
assign MEM[5352] = MEM[4969] + MEM[5050];
assign MEM[5353] = MEM[4970] + MEM[5022];
assign MEM[5354] = MEM[4973] + MEM[5046];
assign MEM[5355] = MEM[4974] + MEM[5071];
assign MEM[5356] = MEM[4981] + MEM[5036];
assign MEM[5357] = MEM[4983] + MEM[5048];
assign MEM[5358] = MEM[4984] + MEM[5030];
assign MEM[5359] = MEM[4985] + MEM[5041];
assign MEM[5360] = MEM[4986] + MEM[5053];
assign MEM[5361] = MEM[4987] + MEM[5029];
assign MEM[5362] = MEM[4991] + MEM[5008];
assign MEM[5363] = MEM[4998] + MEM[5104];
assign MEM[5364] = MEM[4999] + MEM[5087];
assign MEM[5365] = MEM[5002] + MEM[5098];
assign MEM[5366] = MEM[5003] + MEM[5079];
assign MEM[5367] = MEM[5005] + MEM[5032];
assign MEM[5368] = MEM[5006] + MEM[5105];
assign MEM[5369] = MEM[5009] + MEM[5056];
assign MEM[5370] = MEM[5014] + MEM[5062];
assign MEM[5371] = MEM[5015] + MEM[5117];
assign MEM[5372] = MEM[5016] + MEM[5058];
assign MEM[5373] = MEM[5017] + MEM[5077];
assign MEM[5374] = MEM[5018] + MEM[5038];
assign MEM[5375] = MEM[5019] + MEM[5066];
assign MEM[5376] = MEM[5021] + MEM[5115];
assign MEM[5377] = MEM[5023] + MEM[5106];
assign MEM[5378] = MEM[5026] + MEM[5063];
assign MEM[5379] = MEM[5028] + MEM[5097];
assign MEM[5380] = MEM[5031] + MEM[5055];
assign MEM[5381] = MEM[5033] + MEM[5051];
assign MEM[5382] = MEM[5037] + MEM[5129];
assign MEM[5383] = MEM[5039] + MEM[5125];
assign MEM[5384] = MEM[5044] + MEM[5145];
assign MEM[5385] = MEM[5045] + MEM[5100];
assign MEM[5386] = MEM[5049] + MEM[5075];
assign MEM[5387] = MEM[5052] + MEM[5092];
assign MEM[5388] = MEM[5054] + MEM[5180];
assign MEM[5389] = MEM[5057] + MEM[5137];
assign MEM[5390] = MEM[5059] + MEM[5107];
assign MEM[5391] = MEM[5060] + MEM[5134];
assign MEM[5392] = MEM[5061] + MEM[5113];
assign MEM[5393] = MEM[5064] + MEM[5122];
assign MEM[5394] = MEM[5065] + MEM[5116];
assign MEM[5395] = MEM[5067] + MEM[5150];
assign MEM[5396] = MEM[5068] + MEM[5148];
assign MEM[5397] = MEM[5069] + MEM[5188];
assign MEM[5398] = MEM[5070] + MEM[5132];
assign MEM[5399] = MEM[5072] + MEM[5186];
assign MEM[5400] = MEM[5073] + MEM[5120];
assign MEM[5401] = MEM[5074] + MEM[5126];
assign MEM[5402] = MEM[5076] + MEM[5123];
assign MEM[5403] = MEM[5078] + MEM[5141];
assign MEM[5404] = MEM[5080] + MEM[5157];
assign MEM[5405] = MEM[5081] + MEM[5169];
assign MEM[5406] = MEM[5082] + MEM[5168];
assign MEM[5407] = MEM[5083] + MEM[5119];
assign MEM[5408] = MEM[5084] + MEM[5147];
assign MEM[5409] = MEM[5085] + MEM[5140];
assign MEM[5410] = MEM[5086] + MEM[5133];
assign MEM[5411] = MEM[5088] + MEM[5156];
assign MEM[5412] = MEM[5089] + MEM[5139];
assign MEM[5413] = MEM[5090] + MEM[5166];
assign MEM[5414] = MEM[5091] + MEM[5162];
assign MEM[5415] = MEM[5093] + MEM[5161];
assign MEM[5416] = MEM[5094] + MEM[5149];
assign MEM[5417] = MEM[5095] + MEM[5138];
assign MEM[5418] = MEM[5096] + MEM[5164];
assign MEM[5419] = MEM[5099] + MEM[5152];
assign MEM[5420] = MEM[5101] + MEM[5135];
assign MEM[5421] = MEM[5102] + MEM[5144];
assign MEM[5422] = MEM[5103] + MEM[5176];
assign MEM[5423] = MEM[5108] + MEM[5146];
assign MEM[5424] = MEM[5109] + MEM[5170];
assign MEM[5425] = MEM[5110] + MEM[5204];
assign MEM[5426] = MEM[5111] + MEM[5250];
assign MEM[5427] = MEM[5112] + MEM[5182];
assign MEM[5428] = MEM[5114] + MEM[5153];
assign MEM[5429] = MEM[5118] + MEM[5173];
assign MEM[5430] = MEM[5121] + MEM[5158];
assign MEM[5431] = MEM[5124] + MEM[5172];
assign MEM[5432] = MEM[5127] + MEM[5177];
assign MEM[5433] = MEM[5128] + MEM[5181];
assign MEM[5434] = MEM[5130] + MEM[5171];
assign MEM[5435] = MEM[5131] + MEM[5209];
assign MEM[5436] = MEM[5136] + MEM[5185];
assign MEM[5437] = MEM[5142] + MEM[5175];
assign MEM[5438] = MEM[5143] + MEM[5219];
assign MEM[5439] = MEM[5151] + MEM[5205];
assign MEM[5440] = MEM[5154] + MEM[5220];
assign MEM[5441] = MEM[5155] + MEM[5196];
assign MEM[5442] = MEM[5159] + MEM[5237];
assign MEM[5443] = MEM[5160] + MEM[5203];
assign MEM[5444] = MEM[5163] + MEM[5208];
assign MEM[5445] = MEM[5165] + MEM[5249];
assign MEM[5446] = MEM[5167] + MEM[5285];
assign MEM[5447] = MEM[5174] + MEM[5228];
assign MEM[5448] = MEM[5178] + MEM[5215];
assign MEM[5449] = MEM[5179] + MEM[5236];
assign MEM[5450] = MEM[5183] + MEM[5240];
assign MEM[5451] = MEM[5184] + MEM[5267];
assign MEM[5452] = MEM[5187] + MEM[5244];
assign MEM[5453] = MEM[5189] + MEM[5268];
assign MEM[5454] = MEM[5190] + MEM[5247];
assign MEM[5455] = MEM[5191] + MEM[5270];
assign MEM[5456] = MEM[5192] + MEM[5261];
assign MEM[5457] = MEM[5193] + MEM[5278];
assign MEM[5458] = MEM[5194] + MEM[5272];
assign MEM[5459] = MEM[5195] + MEM[5290];
assign MEM[5460] = MEM[5197] + MEM[5287];
assign MEM[5461] = MEM[5198] + MEM[5259];
assign MEM[5462] = MEM[5199] + MEM[5248];
assign MEM[5463] = MEM[5200] + MEM[5264];
assign MEM[5464] = MEM[5201] + MEM[5269];
assign MEM[5465] = MEM[5202] + MEM[5282];
assign MEM[5466] = MEM[5206] + MEM[5262];
assign MEM[5467] = MEM[5207] + MEM[5260];
assign MEM[5468] = MEM[5210] + MEM[5258];
assign MEM[5469] = MEM[5211] + MEM[5307];
assign MEM[5470] = MEM[5212] + MEM[5284];
assign MEM[5471] = MEM[5213] + MEM[5243];
assign MEM[5472] = MEM[5214] + MEM[5273];
assign MEM[5473] = MEM[5216] + MEM[5239];
assign MEM[5474] = MEM[5217] + MEM[5252];
assign MEM[5475] = MEM[5218] + MEM[5253];
assign MEM[5476] = MEM[5221] + MEM[5281];
assign MEM[5477] = MEM[5222] + MEM[5296];
assign MEM[5478] = MEM[5223] + MEM[5279];
assign MEM[5479] = MEM[5224] + MEM[5277];
assign MEM[5480] = MEM[5225] + MEM[5300];
assign MEM[5481] = MEM[5226] + MEM[5256];
assign MEM[5482] = MEM[5227] + MEM[5293];
assign MEM[5483] = MEM[5229] + MEM[5292];
assign MEM[5484] = MEM[5230] + MEM[5298];
assign MEM[5485] = MEM[5231] + MEM[5289];
assign MEM[5486] = MEM[5232] + MEM[5280];
assign MEM[5487] = MEM[5233] + MEM[5303];
assign MEM[5488] = MEM[5234] + MEM[5302];
assign MEM[5489] = MEM[5235] + MEM[5286];
assign MEM[5490] = MEM[5238] + MEM[5291];
assign MEM[5491] = MEM[5241] + MEM[5322];
assign MEM[5492] = MEM[5242] + MEM[5288];
assign MEM[5493] = MEM[5245] + MEM[5310];
assign MEM[5494] = MEM[5246] + MEM[5294];
assign MEM[5495] = MEM[5251] + MEM[5306];
assign MEM[5496] = MEM[5254] + MEM[5301];
assign MEM[5497] = MEM[5255] + MEM[5319];
assign MEM[5498] = MEM[5257] + MEM[5299];
assign MEM[5499] = MEM[5263] + MEM[5317];
assign MEM[5500] = MEM[5265] + MEM[5374];
assign MEM[5501] = MEM[5266] + MEM[5314];
assign MEM[5502] = MEM[5271] + MEM[5309];
assign MEM[5503] = MEM[5274] + MEM[5333];
assign MEM[5504] = MEM[5275] + MEM[5327];
assign MEM[5505] = MEM[5276] + MEM[5324];
assign MEM[5506] = MEM[5283] + MEM[5335];
assign MEM[5507] = MEM[5295] + MEM[5371];
assign MEM[5508] = MEM[5297] + MEM[5403];
assign MEM[5509] = MEM[5304] + MEM[5362];
assign MEM[5510] = MEM[5305] + MEM[5385];
assign MEM[5511] = MEM[5308] + MEM[5368];
assign MEM[5512] = MEM[5311] + MEM[5393];
assign MEM[5513] = MEM[5312] + MEM[5412];
assign MEM[5514] = MEM[5313] + MEM[5400];
assign MEM[5515] = MEM[5315] + MEM[5408];
assign MEM[5516] = MEM[5316] + MEM[5375];
assign MEM[5517] = MEM[5318] + MEM[5365];
assign MEM[5518] = MEM[5320] + MEM[5434];
assign MEM[5519] = MEM[5321] + MEM[5395];
assign MEM[5520] = MEM[5323] + MEM[5382];
assign MEM[5521] = MEM[5325] + MEM[5388];
assign MEM[5522] = MEM[5326] + MEM[5433];
assign MEM[5523] = MEM[5328] + MEM[5384];
assign MEM[5524] = MEM[5329] + MEM[5377];
assign MEM[5525] = MEM[5330] + MEM[5376];
assign MEM[5526] = MEM[5331] + MEM[5396];
assign MEM[5527] = MEM[5332] + MEM[5383];
assign MEM[5528] = MEM[5334] + MEM[5402];
assign MEM[5529] = MEM[5336] + MEM[5390];
assign MEM[5530] = MEM[5337] + MEM[5389];
assign MEM[5531] = MEM[5338] + MEM[5405];
assign MEM[5532] = MEM[5339] + MEM[5404];
assign MEM[5533] = MEM[5340] + MEM[5423];
assign MEM[5534] = MEM[5341] + MEM[5399];
assign MEM[5535] = MEM[5342] + MEM[5378];
assign MEM[5536] = MEM[5343] + MEM[5417];
assign MEM[5537] = MEM[5344] + MEM[5419];
assign MEM[5538] = MEM[5345] + MEM[5411];
assign MEM[5539] = MEM[5346] + MEM[5392];
assign MEM[5540] = MEM[5347] + MEM[5397];
assign MEM[5541] = MEM[5348] + MEM[5406];
assign MEM[5542] = MEM[5349] + MEM[5394];
assign MEM[5543] = MEM[5350] + MEM[5421];
assign MEM[5544] = MEM[5351] + MEM[5414];
assign MEM[5545] = MEM[5352] + MEM[5428];
assign MEM[5546] = MEM[5353] + MEM[5413];
assign MEM[5547] = MEM[5354] + MEM[5416];
assign MEM[5548] = MEM[5355] + MEM[5437];
assign MEM[5549] = MEM[5356] + MEM[5398];
assign MEM[5550] = MEM[5357] + MEM[5418];
assign MEM[5551] = MEM[5358] + MEM[5415];
assign MEM[5552] = MEM[5359] + MEM[5409];
assign MEM[5553] = MEM[5360] + MEM[5429];
assign MEM[5554] = MEM[5361] + MEM[5401];
assign MEM[5555] = MEM[5363] + MEM[5439];
assign MEM[5556] = MEM[5364] + MEM[5444];
assign MEM[5557] = MEM[5366] + MEM[5430];
assign MEM[5558] = MEM[5367] + MEM[5410];
assign MEM[5559] = MEM[5369] + MEM[5424];
assign MEM[5560] = MEM[5370] + MEM[5431];
assign MEM[5561] = MEM[5372] + MEM[5427];
assign MEM[5562] = MEM[5373] + MEM[5436];
assign MEM[5563] = MEM[5379] + MEM[5438];
assign MEM[5564] = MEM[5380] + MEM[5425];
assign MEM[5565] = MEM[5381] + MEM[5422];
assign MEM[5566] = MEM[5386] + MEM[5432];
assign MEM[5567] = MEM[5387] + MEM[5441];
assign MEM[5568] = MEM[5391] + MEM[5449];
assign MEM[5569] = MEM[5407] + MEM[5440];
assign MEM[5570] = MEM[5420] + MEM[5447];
assign MEM[5571] = MEM[5426] + MEM[5516];
assign MEM[5572] = MEM[5435] + MEM[5509];
assign MEM[5573] = MEM[5442] + MEM[5511];
assign MEM[5574] = MEM[5443] + MEM[5507];
assign MEM[5575] = MEM[5445] + MEM[5535];
assign MEM[5576] = MEM[5446] + MEM[5527];
assign MEM[5577] = MEM[5448] + MEM[5514];
assign MEM[5578] = MEM[5450] + MEM[5539];
assign MEM[5579] = MEM[5451] + MEM[5528];
assign MEM[5580] = MEM[5452] + MEM[5517];
assign MEM[5581] = MEM[5453] + MEM[5524];
assign MEM[5582] = MEM[5454] + MEM[5510];
assign MEM[5583] = MEM[5455] + MEM[5519];
assign MEM[5584] = MEM[5456] + MEM[5532];
assign MEM[5585] = MEM[5457] + MEM[5525];
assign MEM[5586] = MEM[5458] + MEM[5538];
assign MEM[5587] = MEM[5459] + MEM[5549];
assign MEM[5588] = MEM[5460] + MEM[5515];
assign MEM[5589] = MEM[5461] + MEM[5513];
assign MEM[5590] = MEM[5462] + MEM[5512];
assign MEM[5591] = MEM[5463] + MEM[5508];
assign MEM[5592] = MEM[5464] + MEM[5542];
assign MEM[5593] = MEM[5465] + MEM[5536];
assign MEM[5594] = MEM[5466] + MEM[5543];
assign MEM[5595] = MEM[5467] + MEM[5547];
assign MEM[5596] = MEM[5468] + MEM[5520];
assign MEM[5597] = MEM[5469] + MEM[5554];
assign MEM[5598] = MEM[5470] + MEM[5544];
assign MEM[5599] = MEM[5471] + MEM[5533];
assign MEM[5600] = MEM[5472] + MEM[5526];
assign MEM[5601] = MEM[5473] + MEM[5523];
assign MEM[5602] = MEM[5474] + MEM[5552];
assign MEM[5603] = MEM[5475] + MEM[5518];
assign MEM[5604] = MEM[5476] + MEM[5560];
assign MEM[5605] = MEM[5477] + MEM[5530];
assign MEM[5606] = MEM[5478] + MEM[5529];
assign MEM[5607] = MEM[5479] + MEM[5521];
assign MEM[5608] = MEM[5480] + MEM[5550];
assign MEM[5609] = MEM[5481] + MEM[5531];
assign MEM[5610] = MEM[5482] + MEM[5553];
assign MEM[5611] = MEM[5483] + MEM[5559];
assign MEM[5612] = MEM[5484] + MEM[5534];
assign MEM[5613] = MEM[5485] + MEM[5541];
assign MEM[5614] = MEM[5486] + MEM[5545];
assign MEM[5615] = MEM[5487] + MEM[5551];
assign MEM[5616] = MEM[5488] + MEM[5555];
assign MEM[5617] = MEM[5489] + MEM[5522];
assign MEM[5618] = MEM[5490] + MEM[5540];
assign MEM[5619] = MEM[5491] + MEM[5567];
assign MEM[5620] = MEM[5492] + MEM[5548];
assign MEM[5621] = MEM[5493] + MEM[5561];
assign MEM[5622] = MEM[5494] + MEM[5546];
assign MEM[5623] = MEM[5495] + MEM[5537];
assign MEM[5624] = MEM[5496] + MEM[5558];
assign MEM[5625] = MEM[5497] + MEM[5566];
assign MEM[5626] = MEM[5498] + MEM[5563];
assign MEM[5627] = MEM[5499] + MEM[5556];
assign MEM[5628] = MEM[5500] + MEM[5569];
assign MEM[5629] = MEM[5501] + MEM[5557];
assign MEM[5630] = MEM[5502] + MEM[5565];
assign MEM[5631] = MEM[5503] + MEM[5570];
assign MEM[5632] = MEM[5504] + MEM[5564];
assign MEM[5633] = MEM[5505] + MEM[5562];
assign MEM[5634] = MEM[5506] + MEM[5568];
assign output_vector[0] = MEM[5611];
assign output_vector[1] = MEM[5602];
assign output_vector[2] = MEM[5618];
assign output_vector[3] = MEM[5603];
assign output_vector[4] = MEM[5597];
assign output_vector[5] = MEM[5576];
assign output_vector[6] = MEM[5595];
assign output_vector[7] = MEM[5580];
assign output_vector[8] = MEM[5617];
assign output_vector[9] = MEM[5616];
assign output_vector[10] = MEM[5599];
assign output_vector[11] = MEM[5627];
assign output_vector[12] = MEM[5575];
assign output_vector[13] = MEM[5613];
assign output_vector[14] = MEM[5571];
assign output_vector[15] = MEM[5623];
assign output_vector[16] = MEM[5600];
assign output_vector[17] = MEM[5584];
assign output_vector[18] = MEM[5588];
assign output_vector[19] = MEM[5631];
assign output_vector[20] = MEM[5589];
assign output_vector[21] = MEM[5620];
assign output_vector[22] = MEM[5582];
assign output_vector[23] = MEM[5590];
assign output_vector[24] = MEM[5621];
assign output_vector[25] = MEM[5610];
assign output_vector[26] = MEM[5614];
assign output_vector[27] = MEM[5594];
assign output_vector[28] = MEM[5573];
assign output_vector[29] = MEM[5578];
assign output_vector[30] = MEM[5591];
assign output_vector[31] = MEM[5629];
assign output_vector[32] = MEM[5633];
assign output_vector[33] = MEM[5607];
assign output_vector[34] = MEM[5609];
assign output_vector[35] = MEM[5572];
assign output_vector[36] = MEM[5615];
assign output_vector[37] = MEM[5632];
assign output_vector[38] = MEM[5628];
assign output_vector[39] = MEM[5596];
assign output_vector[40] = MEM[5622];
assign output_vector[41] = MEM[5583];
assign output_vector[42] = MEM[5574];
assign output_vector[43] = MEM[5601];
assign output_vector[44] = MEM[5586];
assign output_vector[45] = MEM[5624];
assign output_vector[46] = MEM[5630];
assign output_vector[47] = MEM[5606];
assign output_vector[48] = MEM[5581];
assign output_vector[49] = MEM[5625];
assign output_vector[50] = MEM[5585];
assign output_vector[51] = MEM[5598];
assign output_vector[52] = MEM[5593];
assign output_vector[53] = MEM[5608];
assign output_vector[54] = MEM[5577];
assign output_vector[55] = MEM[5634];
assign output_vector[56] = MEM[5579];
assign output_vector[57] = MEM[5587];
assign output_vector[58] = MEM[5605];
assign output_vector[59] = MEM[5619];
assign output_vector[60] = MEM[5626];
assign output_vector[61] = MEM[5592];
assign output_vector[62] = MEM[5604];
assign output_vector[63] = MEM[5612];

endmodule
