// Verilog module
module matrix_mult_optimized_64x784_8_49770#(
    parameter ROWS = 64,
    parameter COLS = 784,
    parameter MEM_SIZE = 49770,
    parameter input_bit_width = 9,
    parameter output_bit_width = 26
)(
    input wire signed [input_bit_width-1:0] input_vector [0: COLS-1],
   output wire signed [output_bit_width-1:0] output_vector [0: ROWS-1]
);

wire signed [output_bit_width-1:0] MEM [0:MEM_SIZE];

assign MEM[0] = -(input_vector[0] << 7);
assign MEM[1] = input_vector[0] << 6;
assign MEM[2] = input_vector[0] << 5;
assign MEM[3] = input_vector[0] << 4;
assign MEM[4] = input_vector[0] << 3;
assign MEM[5] = input_vector[0] << 2;
assign MEM[6] = input_vector[0] << 1;
assign MEM[7] = input_vector[0] << 0;
assign MEM[8] = -(input_vector[1] << 7);
assign MEM[9] = input_vector[1] << 6;
assign MEM[10] = input_vector[1] << 5;
assign MEM[11] = input_vector[1] << 4;
assign MEM[12] = input_vector[1] << 3;
assign MEM[13] = input_vector[1] << 2;
assign MEM[14] = input_vector[1] << 1;
assign MEM[15] = input_vector[1] << 0;
assign MEM[16] = -(input_vector[2] << 7);
assign MEM[17] = input_vector[2] << 6;
assign MEM[18] = input_vector[2] << 5;
assign MEM[19] = input_vector[2] << 4;
assign MEM[20] = input_vector[2] << 3;
assign MEM[21] = input_vector[2] << 2;
assign MEM[22] = input_vector[2] << 1;
assign MEM[23] = input_vector[2] << 0;
assign MEM[24] = -(input_vector[3] << 7);
assign MEM[25] = input_vector[3] << 6;
assign MEM[26] = input_vector[3] << 5;
assign MEM[27] = input_vector[3] << 4;
assign MEM[28] = input_vector[3] << 3;
assign MEM[29] = input_vector[3] << 2;
assign MEM[30] = input_vector[3] << 1;
assign MEM[31] = input_vector[3] << 0;
assign MEM[32] = -(input_vector[4] << 7);
assign MEM[33] = input_vector[4] << 6;
assign MEM[34] = input_vector[4] << 5;
assign MEM[35] = input_vector[4] << 4;
assign MEM[36] = input_vector[4] << 3;
assign MEM[37] = input_vector[4] << 2;
assign MEM[38] = input_vector[4] << 1;
assign MEM[39] = input_vector[4] << 0;
assign MEM[40] = -(input_vector[5] << 7);
assign MEM[41] = input_vector[5] << 6;
assign MEM[42] = input_vector[5] << 5;
assign MEM[43] = input_vector[5] << 4;
assign MEM[44] = input_vector[5] << 3;
assign MEM[45] = input_vector[5] << 2;
assign MEM[46] = input_vector[5] << 1;
assign MEM[47] = input_vector[5] << 0;
assign MEM[48] = -(input_vector[6] << 7);
assign MEM[49] = input_vector[6] << 6;
assign MEM[50] = input_vector[6] << 5;
assign MEM[51] = input_vector[6] << 4;
assign MEM[52] = input_vector[6] << 3;
assign MEM[53] = input_vector[6] << 2;
assign MEM[54] = input_vector[6] << 1;
assign MEM[55] = input_vector[6] << 0;
assign MEM[56] = -(input_vector[7] << 7);
assign MEM[57] = input_vector[7] << 6;
assign MEM[58] = input_vector[7] << 5;
assign MEM[59] = input_vector[7] << 4;
assign MEM[60] = input_vector[7] << 3;
assign MEM[61] = input_vector[7] << 2;
assign MEM[62] = input_vector[7] << 1;
assign MEM[63] = input_vector[7] << 0;
assign MEM[64] = -(input_vector[8] << 7);
assign MEM[65] = input_vector[8] << 6;
assign MEM[66] = input_vector[8] << 5;
assign MEM[67] = input_vector[8] << 4;
assign MEM[68] = input_vector[8] << 3;
assign MEM[69] = input_vector[8] << 2;
assign MEM[70] = input_vector[8] << 1;
assign MEM[71] = input_vector[8] << 0;
assign MEM[72] = -(input_vector[9] << 7);
assign MEM[73] = input_vector[9] << 6;
assign MEM[74] = input_vector[9] << 5;
assign MEM[75] = input_vector[9] << 4;
assign MEM[76] = input_vector[9] << 3;
assign MEM[77] = input_vector[9] << 2;
assign MEM[78] = input_vector[9] << 1;
assign MEM[79] = input_vector[9] << 0;
assign MEM[80] = -(input_vector[10] << 7);
assign MEM[81] = input_vector[10] << 6;
assign MEM[82] = input_vector[10] << 5;
assign MEM[83] = input_vector[10] << 4;
assign MEM[84] = input_vector[10] << 3;
assign MEM[85] = input_vector[10] << 2;
assign MEM[86] = input_vector[10] << 1;
assign MEM[87] = input_vector[10] << 0;
assign MEM[88] = -(input_vector[11] << 7);
assign MEM[89] = input_vector[11] << 6;
assign MEM[90] = input_vector[11] << 5;
assign MEM[91] = input_vector[11] << 4;
assign MEM[92] = input_vector[11] << 3;
assign MEM[93] = input_vector[11] << 2;
assign MEM[94] = input_vector[11] << 1;
assign MEM[95] = input_vector[11] << 0;
assign MEM[96] = -(input_vector[12] << 7);
assign MEM[97] = input_vector[12] << 6;
assign MEM[98] = input_vector[12] << 5;
assign MEM[99] = input_vector[12] << 4;
assign MEM[100] = input_vector[12] << 3;
assign MEM[101] = input_vector[12] << 2;
assign MEM[102] = input_vector[12] << 1;
assign MEM[103] = input_vector[12] << 0;
assign MEM[104] = -(input_vector[13] << 7);
assign MEM[105] = input_vector[13] << 6;
assign MEM[106] = input_vector[13] << 5;
assign MEM[107] = input_vector[13] << 4;
assign MEM[108] = input_vector[13] << 3;
assign MEM[109] = input_vector[13] << 2;
assign MEM[110] = input_vector[13] << 1;
assign MEM[111] = input_vector[13] << 0;
assign MEM[112] = -(input_vector[14] << 7);
assign MEM[113] = input_vector[14] << 6;
assign MEM[114] = input_vector[14] << 5;
assign MEM[115] = input_vector[14] << 4;
assign MEM[116] = input_vector[14] << 3;
assign MEM[117] = input_vector[14] << 2;
assign MEM[118] = input_vector[14] << 1;
assign MEM[119] = input_vector[14] << 0;
assign MEM[120] = -(input_vector[15] << 7);
assign MEM[121] = input_vector[15] << 6;
assign MEM[122] = input_vector[15] << 5;
assign MEM[123] = input_vector[15] << 4;
assign MEM[124] = input_vector[15] << 3;
assign MEM[125] = input_vector[15] << 2;
assign MEM[126] = input_vector[15] << 1;
assign MEM[127] = input_vector[15] << 0;
assign MEM[128] = -(input_vector[16] << 7);
assign MEM[129] = input_vector[16] << 6;
assign MEM[130] = input_vector[16] << 5;
assign MEM[131] = input_vector[16] << 4;
assign MEM[132] = input_vector[16] << 3;
assign MEM[133] = input_vector[16] << 2;
assign MEM[134] = input_vector[16] << 1;
assign MEM[135] = input_vector[16] << 0;
assign MEM[136] = -(input_vector[17] << 7);
assign MEM[137] = input_vector[17] << 6;
assign MEM[138] = input_vector[17] << 5;
assign MEM[139] = input_vector[17] << 4;
assign MEM[140] = input_vector[17] << 3;
assign MEM[141] = input_vector[17] << 2;
assign MEM[142] = input_vector[17] << 1;
assign MEM[143] = input_vector[17] << 0;
assign MEM[144] = -(input_vector[18] << 7);
assign MEM[145] = input_vector[18] << 6;
assign MEM[146] = input_vector[18] << 5;
assign MEM[147] = input_vector[18] << 4;
assign MEM[148] = input_vector[18] << 3;
assign MEM[149] = input_vector[18] << 2;
assign MEM[150] = input_vector[18] << 1;
assign MEM[151] = input_vector[18] << 0;
assign MEM[152] = -(input_vector[19] << 7);
assign MEM[153] = input_vector[19] << 6;
assign MEM[154] = input_vector[19] << 5;
assign MEM[155] = input_vector[19] << 4;
assign MEM[156] = input_vector[19] << 3;
assign MEM[157] = input_vector[19] << 2;
assign MEM[158] = input_vector[19] << 1;
assign MEM[159] = input_vector[19] << 0;
assign MEM[160] = -(input_vector[20] << 7);
assign MEM[161] = input_vector[20] << 6;
assign MEM[162] = input_vector[20] << 5;
assign MEM[163] = input_vector[20] << 4;
assign MEM[164] = input_vector[20] << 3;
assign MEM[165] = input_vector[20] << 2;
assign MEM[166] = input_vector[20] << 1;
assign MEM[167] = input_vector[20] << 0;
assign MEM[168] = -(input_vector[21] << 7);
assign MEM[169] = input_vector[21] << 6;
assign MEM[170] = input_vector[21] << 5;
assign MEM[171] = input_vector[21] << 4;
assign MEM[172] = input_vector[21] << 3;
assign MEM[173] = input_vector[21] << 2;
assign MEM[174] = input_vector[21] << 1;
assign MEM[175] = input_vector[21] << 0;
assign MEM[176] = -(input_vector[22] << 7);
assign MEM[177] = input_vector[22] << 6;
assign MEM[178] = input_vector[22] << 5;
assign MEM[179] = input_vector[22] << 4;
assign MEM[180] = input_vector[22] << 3;
assign MEM[181] = input_vector[22] << 2;
assign MEM[182] = input_vector[22] << 1;
assign MEM[183] = input_vector[22] << 0;
assign MEM[184] = -(input_vector[23] << 7);
assign MEM[185] = input_vector[23] << 6;
assign MEM[186] = input_vector[23] << 5;
assign MEM[187] = input_vector[23] << 4;
assign MEM[188] = input_vector[23] << 3;
assign MEM[189] = input_vector[23] << 2;
assign MEM[190] = input_vector[23] << 1;
assign MEM[191] = input_vector[23] << 0;
assign MEM[192] = -(input_vector[24] << 7);
assign MEM[193] = input_vector[24] << 6;
assign MEM[194] = input_vector[24] << 5;
assign MEM[195] = input_vector[24] << 4;
assign MEM[196] = input_vector[24] << 3;
assign MEM[197] = input_vector[24] << 2;
assign MEM[198] = input_vector[24] << 1;
assign MEM[199] = input_vector[24] << 0;
assign MEM[200] = -(input_vector[25] << 7);
assign MEM[201] = input_vector[25] << 6;
assign MEM[202] = input_vector[25] << 5;
assign MEM[203] = input_vector[25] << 4;
assign MEM[204] = input_vector[25] << 3;
assign MEM[205] = input_vector[25] << 2;
assign MEM[206] = input_vector[25] << 1;
assign MEM[207] = input_vector[25] << 0;
assign MEM[208] = -(input_vector[26] << 7);
assign MEM[209] = input_vector[26] << 6;
assign MEM[210] = input_vector[26] << 5;
assign MEM[211] = input_vector[26] << 4;
assign MEM[212] = input_vector[26] << 3;
assign MEM[213] = input_vector[26] << 2;
assign MEM[214] = input_vector[26] << 1;
assign MEM[215] = input_vector[26] << 0;
assign MEM[216] = -(input_vector[27] << 7);
assign MEM[217] = input_vector[27] << 6;
assign MEM[218] = input_vector[27] << 5;
assign MEM[219] = input_vector[27] << 4;
assign MEM[220] = input_vector[27] << 3;
assign MEM[221] = input_vector[27] << 2;
assign MEM[222] = input_vector[27] << 1;
assign MEM[223] = input_vector[27] << 0;
assign MEM[224] = -(input_vector[28] << 7);
assign MEM[225] = input_vector[28] << 6;
assign MEM[226] = input_vector[28] << 5;
assign MEM[227] = input_vector[28] << 4;
assign MEM[228] = input_vector[28] << 3;
assign MEM[229] = input_vector[28] << 2;
assign MEM[230] = input_vector[28] << 1;
assign MEM[231] = input_vector[28] << 0;
assign MEM[232] = -(input_vector[29] << 7);
assign MEM[233] = input_vector[29] << 6;
assign MEM[234] = input_vector[29] << 5;
assign MEM[235] = input_vector[29] << 4;
assign MEM[236] = input_vector[29] << 3;
assign MEM[237] = input_vector[29] << 2;
assign MEM[238] = input_vector[29] << 1;
assign MEM[239] = input_vector[29] << 0;
assign MEM[240] = -(input_vector[30] << 7);
assign MEM[241] = input_vector[30] << 6;
assign MEM[242] = input_vector[30] << 5;
assign MEM[243] = input_vector[30] << 4;
assign MEM[244] = input_vector[30] << 3;
assign MEM[245] = input_vector[30] << 2;
assign MEM[246] = input_vector[30] << 1;
assign MEM[247] = input_vector[30] << 0;
assign MEM[248] = -(input_vector[31] << 7);
assign MEM[249] = input_vector[31] << 6;
assign MEM[250] = input_vector[31] << 5;
assign MEM[251] = input_vector[31] << 4;
assign MEM[252] = input_vector[31] << 3;
assign MEM[253] = input_vector[31] << 2;
assign MEM[254] = input_vector[31] << 1;
assign MEM[255] = input_vector[31] << 0;
assign MEM[256] = -(input_vector[32] << 7);
assign MEM[257] = input_vector[32] << 6;
assign MEM[258] = input_vector[32] << 5;
assign MEM[259] = input_vector[32] << 4;
assign MEM[260] = input_vector[32] << 3;
assign MEM[261] = input_vector[32] << 2;
assign MEM[262] = input_vector[32] << 1;
assign MEM[263] = input_vector[32] << 0;
assign MEM[264] = -(input_vector[33] << 7);
assign MEM[265] = input_vector[33] << 6;
assign MEM[266] = input_vector[33] << 5;
assign MEM[267] = input_vector[33] << 4;
assign MEM[268] = input_vector[33] << 3;
assign MEM[269] = input_vector[33] << 2;
assign MEM[270] = input_vector[33] << 1;
assign MEM[271] = input_vector[33] << 0;
assign MEM[272] = -(input_vector[34] << 7);
assign MEM[273] = input_vector[34] << 6;
assign MEM[274] = input_vector[34] << 5;
assign MEM[275] = input_vector[34] << 4;
assign MEM[276] = input_vector[34] << 3;
assign MEM[277] = input_vector[34] << 2;
assign MEM[278] = input_vector[34] << 1;
assign MEM[279] = input_vector[34] << 0;
assign MEM[280] = -(input_vector[35] << 7);
assign MEM[281] = input_vector[35] << 6;
assign MEM[282] = input_vector[35] << 5;
assign MEM[283] = input_vector[35] << 4;
assign MEM[284] = input_vector[35] << 3;
assign MEM[285] = input_vector[35] << 2;
assign MEM[286] = input_vector[35] << 1;
assign MEM[287] = input_vector[35] << 0;
assign MEM[288] = -(input_vector[36] << 7);
assign MEM[289] = input_vector[36] << 6;
assign MEM[290] = input_vector[36] << 5;
assign MEM[291] = input_vector[36] << 4;
assign MEM[292] = input_vector[36] << 3;
assign MEM[293] = input_vector[36] << 2;
assign MEM[294] = input_vector[36] << 1;
assign MEM[295] = input_vector[36] << 0;
assign MEM[296] = -(input_vector[37] << 7);
assign MEM[297] = input_vector[37] << 6;
assign MEM[298] = input_vector[37] << 5;
assign MEM[299] = input_vector[37] << 4;
assign MEM[300] = input_vector[37] << 3;
assign MEM[301] = input_vector[37] << 2;
assign MEM[302] = input_vector[37] << 1;
assign MEM[303] = input_vector[37] << 0;
assign MEM[304] = -(input_vector[38] << 7);
assign MEM[305] = input_vector[38] << 6;
assign MEM[306] = input_vector[38] << 5;
assign MEM[307] = input_vector[38] << 4;
assign MEM[308] = input_vector[38] << 3;
assign MEM[309] = input_vector[38] << 2;
assign MEM[310] = input_vector[38] << 1;
assign MEM[311] = input_vector[38] << 0;
assign MEM[312] = -(input_vector[39] << 7);
assign MEM[313] = input_vector[39] << 6;
assign MEM[314] = input_vector[39] << 5;
assign MEM[315] = input_vector[39] << 4;
assign MEM[316] = input_vector[39] << 3;
assign MEM[317] = input_vector[39] << 2;
assign MEM[318] = input_vector[39] << 1;
assign MEM[319] = input_vector[39] << 0;
assign MEM[320] = -(input_vector[40] << 7);
assign MEM[321] = input_vector[40] << 6;
assign MEM[322] = input_vector[40] << 5;
assign MEM[323] = input_vector[40] << 4;
assign MEM[324] = input_vector[40] << 3;
assign MEM[325] = input_vector[40] << 2;
assign MEM[326] = input_vector[40] << 1;
assign MEM[327] = input_vector[40] << 0;
assign MEM[328] = -(input_vector[41] << 7);
assign MEM[329] = input_vector[41] << 6;
assign MEM[330] = input_vector[41] << 5;
assign MEM[331] = input_vector[41] << 4;
assign MEM[332] = input_vector[41] << 3;
assign MEM[333] = input_vector[41] << 2;
assign MEM[334] = input_vector[41] << 1;
assign MEM[335] = input_vector[41] << 0;
assign MEM[336] = -(input_vector[42] << 7);
assign MEM[337] = input_vector[42] << 6;
assign MEM[338] = input_vector[42] << 5;
assign MEM[339] = input_vector[42] << 4;
assign MEM[340] = input_vector[42] << 3;
assign MEM[341] = input_vector[42] << 2;
assign MEM[342] = input_vector[42] << 1;
assign MEM[343] = input_vector[42] << 0;
assign MEM[344] = -(input_vector[43] << 7);
assign MEM[345] = input_vector[43] << 6;
assign MEM[346] = input_vector[43] << 5;
assign MEM[347] = input_vector[43] << 4;
assign MEM[348] = input_vector[43] << 3;
assign MEM[349] = input_vector[43] << 2;
assign MEM[350] = input_vector[43] << 1;
assign MEM[351] = input_vector[43] << 0;
assign MEM[352] = -(input_vector[44] << 7);
assign MEM[353] = input_vector[44] << 6;
assign MEM[354] = input_vector[44] << 5;
assign MEM[355] = input_vector[44] << 4;
assign MEM[356] = input_vector[44] << 3;
assign MEM[357] = input_vector[44] << 2;
assign MEM[358] = input_vector[44] << 1;
assign MEM[359] = input_vector[44] << 0;
assign MEM[360] = -(input_vector[45] << 7);
assign MEM[361] = input_vector[45] << 6;
assign MEM[362] = input_vector[45] << 5;
assign MEM[363] = input_vector[45] << 4;
assign MEM[364] = input_vector[45] << 3;
assign MEM[365] = input_vector[45] << 2;
assign MEM[366] = input_vector[45] << 1;
assign MEM[367] = input_vector[45] << 0;
assign MEM[368] = -(input_vector[46] << 7);
assign MEM[369] = input_vector[46] << 6;
assign MEM[370] = input_vector[46] << 5;
assign MEM[371] = input_vector[46] << 4;
assign MEM[372] = input_vector[46] << 3;
assign MEM[373] = input_vector[46] << 2;
assign MEM[374] = input_vector[46] << 1;
assign MEM[375] = input_vector[46] << 0;
assign MEM[376] = -(input_vector[47] << 7);
assign MEM[377] = input_vector[47] << 6;
assign MEM[378] = input_vector[47] << 5;
assign MEM[379] = input_vector[47] << 4;
assign MEM[380] = input_vector[47] << 3;
assign MEM[381] = input_vector[47] << 2;
assign MEM[382] = input_vector[47] << 1;
assign MEM[383] = input_vector[47] << 0;
assign MEM[384] = -(input_vector[48] << 7);
assign MEM[385] = input_vector[48] << 6;
assign MEM[386] = input_vector[48] << 5;
assign MEM[387] = input_vector[48] << 4;
assign MEM[388] = input_vector[48] << 3;
assign MEM[389] = input_vector[48] << 2;
assign MEM[390] = input_vector[48] << 1;
assign MEM[391] = input_vector[48] << 0;
assign MEM[392] = -(input_vector[49] << 7);
assign MEM[393] = input_vector[49] << 6;
assign MEM[394] = input_vector[49] << 5;
assign MEM[395] = input_vector[49] << 4;
assign MEM[396] = input_vector[49] << 3;
assign MEM[397] = input_vector[49] << 2;
assign MEM[398] = input_vector[49] << 1;
assign MEM[399] = input_vector[49] << 0;
assign MEM[400] = -(input_vector[50] << 7);
assign MEM[401] = input_vector[50] << 6;
assign MEM[402] = input_vector[50] << 5;
assign MEM[403] = input_vector[50] << 4;
assign MEM[404] = input_vector[50] << 3;
assign MEM[405] = input_vector[50] << 2;
assign MEM[406] = input_vector[50] << 1;
assign MEM[407] = input_vector[50] << 0;
assign MEM[408] = -(input_vector[51] << 7);
assign MEM[409] = input_vector[51] << 6;
assign MEM[410] = input_vector[51] << 5;
assign MEM[411] = input_vector[51] << 4;
assign MEM[412] = input_vector[51] << 3;
assign MEM[413] = input_vector[51] << 2;
assign MEM[414] = input_vector[51] << 1;
assign MEM[415] = input_vector[51] << 0;
assign MEM[416] = -(input_vector[52] << 7);
assign MEM[417] = input_vector[52] << 6;
assign MEM[418] = input_vector[52] << 5;
assign MEM[419] = input_vector[52] << 4;
assign MEM[420] = input_vector[52] << 3;
assign MEM[421] = input_vector[52] << 2;
assign MEM[422] = input_vector[52] << 1;
assign MEM[423] = input_vector[52] << 0;
assign MEM[424] = -(input_vector[53] << 7);
assign MEM[425] = input_vector[53] << 6;
assign MEM[426] = input_vector[53] << 5;
assign MEM[427] = input_vector[53] << 4;
assign MEM[428] = input_vector[53] << 3;
assign MEM[429] = input_vector[53] << 2;
assign MEM[430] = input_vector[53] << 1;
assign MEM[431] = input_vector[53] << 0;
assign MEM[432] = -(input_vector[54] << 7);
assign MEM[433] = input_vector[54] << 6;
assign MEM[434] = input_vector[54] << 5;
assign MEM[435] = input_vector[54] << 4;
assign MEM[436] = input_vector[54] << 3;
assign MEM[437] = input_vector[54] << 2;
assign MEM[438] = input_vector[54] << 1;
assign MEM[439] = input_vector[54] << 0;
assign MEM[440] = -(input_vector[55] << 7);
assign MEM[441] = input_vector[55] << 6;
assign MEM[442] = input_vector[55] << 5;
assign MEM[443] = input_vector[55] << 4;
assign MEM[444] = input_vector[55] << 3;
assign MEM[445] = input_vector[55] << 2;
assign MEM[446] = input_vector[55] << 1;
assign MEM[447] = input_vector[55] << 0;
assign MEM[448] = -(input_vector[56] << 7);
assign MEM[449] = input_vector[56] << 6;
assign MEM[450] = input_vector[56] << 5;
assign MEM[451] = input_vector[56] << 4;
assign MEM[452] = input_vector[56] << 3;
assign MEM[453] = input_vector[56] << 2;
assign MEM[454] = input_vector[56] << 1;
assign MEM[455] = input_vector[56] << 0;
assign MEM[456] = -(input_vector[57] << 7);
assign MEM[457] = input_vector[57] << 6;
assign MEM[458] = input_vector[57] << 5;
assign MEM[459] = input_vector[57] << 4;
assign MEM[460] = input_vector[57] << 3;
assign MEM[461] = input_vector[57] << 2;
assign MEM[462] = input_vector[57] << 1;
assign MEM[463] = input_vector[57] << 0;
assign MEM[464] = -(input_vector[58] << 7);
assign MEM[465] = input_vector[58] << 6;
assign MEM[466] = input_vector[58] << 5;
assign MEM[467] = input_vector[58] << 4;
assign MEM[468] = input_vector[58] << 3;
assign MEM[469] = input_vector[58] << 2;
assign MEM[470] = input_vector[58] << 1;
assign MEM[471] = input_vector[58] << 0;
assign MEM[472] = -(input_vector[59] << 7);
assign MEM[473] = input_vector[59] << 6;
assign MEM[474] = input_vector[59] << 5;
assign MEM[475] = input_vector[59] << 4;
assign MEM[476] = input_vector[59] << 3;
assign MEM[477] = input_vector[59] << 2;
assign MEM[478] = input_vector[59] << 1;
assign MEM[479] = input_vector[59] << 0;
assign MEM[480] = -(input_vector[60] << 7);
assign MEM[481] = input_vector[60] << 6;
assign MEM[482] = input_vector[60] << 5;
assign MEM[483] = input_vector[60] << 4;
assign MEM[484] = input_vector[60] << 3;
assign MEM[485] = input_vector[60] << 2;
assign MEM[486] = input_vector[60] << 1;
assign MEM[487] = input_vector[60] << 0;
assign MEM[488] = -(input_vector[61] << 7);
assign MEM[489] = input_vector[61] << 6;
assign MEM[490] = input_vector[61] << 5;
assign MEM[491] = input_vector[61] << 4;
assign MEM[492] = input_vector[61] << 3;
assign MEM[493] = input_vector[61] << 2;
assign MEM[494] = input_vector[61] << 1;
assign MEM[495] = input_vector[61] << 0;
assign MEM[496] = -(input_vector[62] << 7);
assign MEM[497] = input_vector[62] << 6;
assign MEM[498] = input_vector[62] << 5;
assign MEM[499] = input_vector[62] << 4;
assign MEM[500] = input_vector[62] << 3;
assign MEM[501] = input_vector[62] << 2;
assign MEM[502] = input_vector[62] << 1;
assign MEM[503] = input_vector[62] << 0;
assign MEM[504] = -(input_vector[63] << 7);
assign MEM[505] = input_vector[63] << 6;
assign MEM[506] = input_vector[63] << 5;
assign MEM[507] = input_vector[63] << 4;
assign MEM[508] = input_vector[63] << 3;
assign MEM[509] = input_vector[63] << 2;
assign MEM[510] = input_vector[63] << 1;
assign MEM[511] = input_vector[63] << 0;
assign MEM[512] = -(input_vector[64] << 7);
assign MEM[513] = input_vector[64] << 6;
assign MEM[514] = input_vector[64] << 5;
assign MEM[515] = input_vector[64] << 4;
assign MEM[516] = input_vector[64] << 3;
assign MEM[517] = input_vector[64] << 2;
assign MEM[518] = input_vector[64] << 1;
assign MEM[519] = input_vector[64] << 0;
assign MEM[520] = -(input_vector[65] << 7);
assign MEM[521] = input_vector[65] << 6;
assign MEM[522] = input_vector[65] << 5;
assign MEM[523] = input_vector[65] << 4;
assign MEM[524] = input_vector[65] << 3;
assign MEM[525] = input_vector[65] << 2;
assign MEM[526] = input_vector[65] << 1;
assign MEM[527] = input_vector[65] << 0;
assign MEM[528] = -(input_vector[66] << 7);
assign MEM[529] = input_vector[66] << 6;
assign MEM[530] = input_vector[66] << 5;
assign MEM[531] = input_vector[66] << 4;
assign MEM[532] = input_vector[66] << 3;
assign MEM[533] = input_vector[66] << 2;
assign MEM[534] = input_vector[66] << 1;
assign MEM[535] = input_vector[66] << 0;
assign MEM[536] = -(input_vector[67] << 7);
assign MEM[537] = input_vector[67] << 6;
assign MEM[538] = input_vector[67] << 5;
assign MEM[539] = input_vector[67] << 4;
assign MEM[540] = input_vector[67] << 3;
assign MEM[541] = input_vector[67] << 2;
assign MEM[542] = input_vector[67] << 1;
assign MEM[543] = input_vector[67] << 0;
assign MEM[544] = -(input_vector[68] << 7);
assign MEM[545] = input_vector[68] << 6;
assign MEM[546] = input_vector[68] << 5;
assign MEM[547] = input_vector[68] << 4;
assign MEM[548] = input_vector[68] << 3;
assign MEM[549] = input_vector[68] << 2;
assign MEM[550] = input_vector[68] << 1;
assign MEM[551] = input_vector[68] << 0;
assign MEM[552] = -(input_vector[69] << 7);
assign MEM[553] = input_vector[69] << 6;
assign MEM[554] = input_vector[69] << 5;
assign MEM[555] = input_vector[69] << 4;
assign MEM[556] = input_vector[69] << 3;
assign MEM[557] = input_vector[69] << 2;
assign MEM[558] = input_vector[69] << 1;
assign MEM[559] = input_vector[69] << 0;
assign MEM[560] = -(input_vector[70] << 7);
assign MEM[561] = input_vector[70] << 6;
assign MEM[562] = input_vector[70] << 5;
assign MEM[563] = input_vector[70] << 4;
assign MEM[564] = input_vector[70] << 3;
assign MEM[565] = input_vector[70] << 2;
assign MEM[566] = input_vector[70] << 1;
assign MEM[567] = input_vector[70] << 0;
assign MEM[568] = -(input_vector[71] << 7);
assign MEM[569] = input_vector[71] << 6;
assign MEM[570] = input_vector[71] << 5;
assign MEM[571] = input_vector[71] << 4;
assign MEM[572] = input_vector[71] << 3;
assign MEM[573] = input_vector[71] << 2;
assign MEM[574] = input_vector[71] << 1;
assign MEM[575] = input_vector[71] << 0;
assign MEM[576] = -(input_vector[72] << 7);
assign MEM[577] = input_vector[72] << 6;
assign MEM[578] = input_vector[72] << 5;
assign MEM[579] = input_vector[72] << 4;
assign MEM[580] = input_vector[72] << 3;
assign MEM[581] = input_vector[72] << 2;
assign MEM[582] = input_vector[72] << 1;
assign MEM[583] = input_vector[72] << 0;
assign MEM[584] = -(input_vector[73] << 7);
assign MEM[585] = input_vector[73] << 6;
assign MEM[586] = input_vector[73] << 5;
assign MEM[587] = input_vector[73] << 4;
assign MEM[588] = input_vector[73] << 3;
assign MEM[589] = input_vector[73] << 2;
assign MEM[590] = input_vector[73] << 1;
assign MEM[591] = input_vector[73] << 0;
assign MEM[592] = -(input_vector[74] << 7);
assign MEM[593] = input_vector[74] << 6;
assign MEM[594] = input_vector[74] << 5;
assign MEM[595] = input_vector[74] << 4;
assign MEM[596] = input_vector[74] << 3;
assign MEM[597] = input_vector[74] << 2;
assign MEM[598] = input_vector[74] << 1;
assign MEM[599] = input_vector[74] << 0;
assign MEM[600] = -(input_vector[75] << 7);
assign MEM[601] = input_vector[75] << 6;
assign MEM[602] = input_vector[75] << 5;
assign MEM[603] = input_vector[75] << 4;
assign MEM[604] = input_vector[75] << 3;
assign MEM[605] = input_vector[75] << 2;
assign MEM[606] = input_vector[75] << 1;
assign MEM[607] = input_vector[75] << 0;
assign MEM[608] = -(input_vector[76] << 7);
assign MEM[609] = input_vector[76] << 6;
assign MEM[610] = input_vector[76] << 5;
assign MEM[611] = input_vector[76] << 4;
assign MEM[612] = input_vector[76] << 3;
assign MEM[613] = input_vector[76] << 2;
assign MEM[614] = input_vector[76] << 1;
assign MEM[615] = input_vector[76] << 0;
assign MEM[616] = -(input_vector[77] << 7);
assign MEM[617] = input_vector[77] << 6;
assign MEM[618] = input_vector[77] << 5;
assign MEM[619] = input_vector[77] << 4;
assign MEM[620] = input_vector[77] << 3;
assign MEM[621] = input_vector[77] << 2;
assign MEM[622] = input_vector[77] << 1;
assign MEM[623] = input_vector[77] << 0;
assign MEM[624] = -(input_vector[78] << 7);
assign MEM[625] = input_vector[78] << 6;
assign MEM[626] = input_vector[78] << 5;
assign MEM[627] = input_vector[78] << 4;
assign MEM[628] = input_vector[78] << 3;
assign MEM[629] = input_vector[78] << 2;
assign MEM[630] = input_vector[78] << 1;
assign MEM[631] = input_vector[78] << 0;
assign MEM[632] = -(input_vector[79] << 7);
assign MEM[633] = input_vector[79] << 6;
assign MEM[634] = input_vector[79] << 5;
assign MEM[635] = input_vector[79] << 4;
assign MEM[636] = input_vector[79] << 3;
assign MEM[637] = input_vector[79] << 2;
assign MEM[638] = input_vector[79] << 1;
assign MEM[639] = input_vector[79] << 0;
assign MEM[640] = -(input_vector[80] << 7);
assign MEM[641] = input_vector[80] << 6;
assign MEM[642] = input_vector[80] << 5;
assign MEM[643] = input_vector[80] << 4;
assign MEM[644] = input_vector[80] << 3;
assign MEM[645] = input_vector[80] << 2;
assign MEM[646] = input_vector[80] << 1;
assign MEM[647] = input_vector[80] << 0;
assign MEM[648] = -(input_vector[81] << 7);
assign MEM[649] = input_vector[81] << 6;
assign MEM[650] = input_vector[81] << 5;
assign MEM[651] = input_vector[81] << 4;
assign MEM[652] = input_vector[81] << 3;
assign MEM[653] = input_vector[81] << 2;
assign MEM[654] = input_vector[81] << 1;
assign MEM[655] = input_vector[81] << 0;
assign MEM[656] = -(input_vector[82] << 7);
assign MEM[657] = input_vector[82] << 6;
assign MEM[658] = input_vector[82] << 5;
assign MEM[659] = input_vector[82] << 4;
assign MEM[660] = input_vector[82] << 3;
assign MEM[661] = input_vector[82] << 2;
assign MEM[662] = input_vector[82] << 1;
assign MEM[663] = input_vector[82] << 0;
assign MEM[664] = -(input_vector[83] << 7);
assign MEM[665] = input_vector[83] << 6;
assign MEM[666] = input_vector[83] << 5;
assign MEM[667] = input_vector[83] << 4;
assign MEM[668] = input_vector[83] << 3;
assign MEM[669] = input_vector[83] << 2;
assign MEM[670] = input_vector[83] << 1;
assign MEM[671] = input_vector[83] << 0;
assign MEM[672] = -(input_vector[84] << 7);
assign MEM[673] = input_vector[84] << 6;
assign MEM[674] = input_vector[84] << 5;
assign MEM[675] = input_vector[84] << 4;
assign MEM[676] = input_vector[84] << 3;
assign MEM[677] = input_vector[84] << 2;
assign MEM[678] = input_vector[84] << 1;
assign MEM[679] = input_vector[84] << 0;
assign MEM[680] = -(input_vector[85] << 7);
assign MEM[681] = input_vector[85] << 6;
assign MEM[682] = input_vector[85] << 5;
assign MEM[683] = input_vector[85] << 4;
assign MEM[684] = input_vector[85] << 3;
assign MEM[685] = input_vector[85] << 2;
assign MEM[686] = input_vector[85] << 1;
assign MEM[687] = input_vector[85] << 0;
assign MEM[688] = -(input_vector[86] << 7);
assign MEM[689] = input_vector[86] << 6;
assign MEM[690] = input_vector[86] << 5;
assign MEM[691] = input_vector[86] << 4;
assign MEM[692] = input_vector[86] << 3;
assign MEM[693] = input_vector[86] << 2;
assign MEM[694] = input_vector[86] << 1;
assign MEM[695] = input_vector[86] << 0;
assign MEM[696] = -(input_vector[87] << 7);
assign MEM[697] = input_vector[87] << 6;
assign MEM[698] = input_vector[87] << 5;
assign MEM[699] = input_vector[87] << 4;
assign MEM[700] = input_vector[87] << 3;
assign MEM[701] = input_vector[87] << 2;
assign MEM[702] = input_vector[87] << 1;
assign MEM[703] = input_vector[87] << 0;
assign MEM[704] = -(input_vector[88] << 7);
assign MEM[705] = input_vector[88] << 6;
assign MEM[706] = input_vector[88] << 5;
assign MEM[707] = input_vector[88] << 4;
assign MEM[708] = input_vector[88] << 3;
assign MEM[709] = input_vector[88] << 2;
assign MEM[710] = input_vector[88] << 1;
assign MEM[711] = input_vector[88] << 0;
assign MEM[712] = -(input_vector[89] << 7);
assign MEM[713] = input_vector[89] << 6;
assign MEM[714] = input_vector[89] << 5;
assign MEM[715] = input_vector[89] << 4;
assign MEM[716] = input_vector[89] << 3;
assign MEM[717] = input_vector[89] << 2;
assign MEM[718] = input_vector[89] << 1;
assign MEM[719] = input_vector[89] << 0;
assign MEM[720] = -(input_vector[90] << 7);
assign MEM[721] = input_vector[90] << 6;
assign MEM[722] = input_vector[90] << 5;
assign MEM[723] = input_vector[90] << 4;
assign MEM[724] = input_vector[90] << 3;
assign MEM[725] = input_vector[90] << 2;
assign MEM[726] = input_vector[90] << 1;
assign MEM[727] = input_vector[90] << 0;
assign MEM[728] = -(input_vector[91] << 7);
assign MEM[729] = input_vector[91] << 6;
assign MEM[730] = input_vector[91] << 5;
assign MEM[731] = input_vector[91] << 4;
assign MEM[732] = input_vector[91] << 3;
assign MEM[733] = input_vector[91] << 2;
assign MEM[734] = input_vector[91] << 1;
assign MEM[735] = input_vector[91] << 0;
assign MEM[736] = -(input_vector[92] << 7);
assign MEM[737] = input_vector[92] << 6;
assign MEM[738] = input_vector[92] << 5;
assign MEM[739] = input_vector[92] << 4;
assign MEM[740] = input_vector[92] << 3;
assign MEM[741] = input_vector[92] << 2;
assign MEM[742] = input_vector[92] << 1;
assign MEM[743] = input_vector[92] << 0;
assign MEM[744] = -(input_vector[93] << 7);
assign MEM[745] = input_vector[93] << 6;
assign MEM[746] = input_vector[93] << 5;
assign MEM[747] = input_vector[93] << 4;
assign MEM[748] = input_vector[93] << 3;
assign MEM[749] = input_vector[93] << 2;
assign MEM[750] = input_vector[93] << 1;
assign MEM[751] = input_vector[93] << 0;
assign MEM[752] = -(input_vector[94] << 7);
assign MEM[753] = input_vector[94] << 6;
assign MEM[754] = input_vector[94] << 5;
assign MEM[755] = input_vector[94] << 4;
assign MEM[756] = input_vector[94] << 3;
assign MEM[757] = input_vector[94] << 2;
assign MEM[758] = input_vector[94] << 1;
assign MEM[759] = input_vector[94] << 0;
assign MEM[760] = -(input_vector[95] << 7);
assign MEM[761] = input_vector[95] << 6;
assign MEM[762] = input_vector[95] << 5;
assign MEM[763] = input_vector[95] << 4;
assign MEM[764] = input_vector[95] << 3;
assign MEM[765] = input_vector[95] << 2;
assign MEM[766] = input_vector[95] << 1;
assign MEM[767] = input_vector[95] << 0;
assign MEM[768] = -(input_vector[96] << 7);
assign MEM[769] = input_vector[96] << 6;
assign MEM[770] = input_vector[96] << 5;
assign MEM[771] = input_vector[96] << 4;
assign MEM[772] = input_vector[96] << 3;
assign MEM[773] = input_vector[96] << 2;
assign MEM[774] = input_vector[96] << 1;
assign MEM[775] = input_vector[96] << 0;
assign MEM[776] = -(input_vector[97] << 7);
assign MEM[777] = input_vector[97] << 6;
assign MEM[778] = input_vector[97] << 5;
assign MEM[779] = input_vector[97] << 4;
assign MEM[780] = input_vector[97] << 3;
assign MEM[781] = input_vector[97] << 2;
assign MEM[782] = input_vector[97] << 1;
assign MEM[783] = input_vector[97] << 0;
assign MEM[784] = -(input_vector[98] << 7);
assign MEM[785] = input_vector[98] << 6;
assign MEM[786] = input_vector[98] << 5;
assign MEM[787] = input_vector[98] << 4;
assign MEM[788] = input_vector[98] << 3;
assign MEM[789] = input_vector[98] << 2;
assign MEM[790] = input_vector[98] << 1;
assign MEM[791] = input_vector[98] << 0;
assign MEM[792] = -(input_vector[99] << 7);
assign MEM[793] = input_vector[99] << 6;
assign MEM[794] = input_vector[99] << 5;
assign MEM[795] = input_vector[99] << 4;
assign MEM[796] = input_vector[99] << 3;
assign MEM[797] = input_vector[99] << 2;
assign MEM[798] = input_vector[99] << 1;
assign MEM[799] = input_vector[99] << 0;
assign MEM[800] = -(input_vector[100] << 7);
assign MEM[801] = input_vector[100] << 6;
assign MEM[802] = input_vector[100] << 5;
assign MEM[803] = input_vector[100] << 4;
assign MEM[804] = input_vector[100] << 3;
assign MEM[805] = input_vector[100] << 2;
assign MEM[806] = input_vector[100] << 1;
assign MEM[807] = input_vector[100] << 0;
assign MEM[808] = -(input_vector[101] << 7);
assign MEM[809] = input_vector[101] << 6;
assign MEM[810] = input_vector[101] << 5;
assign MEM[811] = input_vector[101] << 4;
assign MEM[812] = input_vector[101] << 3;
assign MEM[813] = input_vector[101] << 2;
assign MEM[814] = input_vector[101] << 1;
assign MEM[815] = input_vector[101] << 0;
assign MEM[816] = -(input_vector[102] << 7);
assign MEM[817] = input_vector[102] << 6;
assign MEM[818] = input_vector[102] << 5;
assign MEM[819] = input_vector[102] << 4;
assign MEM[820] = input_vector[102] << 3;
assign MEM[821] = input_vector[102] << 2;
assign MEM[822] = input_vector[102] << 1;
assign MEM[823] = input_vector[102] << 0;
assign MEM[824] = -(input_vector[103] << 7);
assign MEM[825] = input_vector[103] << 6;
assign MEM[826] = input_vector[103] << 5;
assign MEM[827] = input_vector[103] << 4;
assign MEM[828] = input_vector[103] << 3;
assign MEM[829] = input_vector[103] << 2;
assign MEM[830] = input_vector[103] << 1;
assign MEM[831] = input_vector[103] << 0;
assign MEM[832] = -(input_vector[104] << 7);
assign MEM[833] = input_vector[104] << 6;
assign MEM[834] = input_vector[104] << 5;
assign MEM[835] = input_vector[104] << 4;
assign MEM[836] = input_vector[104] << 3;
assign MEM[837] = input_vector[104] << 2;
assign MEM[838] = input_vector[104] << 1;
assign MEM[839] = input_vector[104] << 0;
assign MEM[840] = -(input_vector[105] << 7);
assign MEM[841] = input_vector[105] << 6;
assign MEM[842] = input_vector[105] << 5;
assign MEM[843] = input_vector[105] << 4;
assign MEM[844] = input_vector[105] << 3;
assign MEM[845] = input_vector[105] << 2;
assign MEM[846] = input_vector[105] << 1;
assign MEM[847] = input_vector[105] << 0;
assign MEM[848] = -(input_vector[106] << 7);
assign MEM[849] = input_vector[106] << 6;
assign MEM[850] = input_vector[106] << 5;
assign MEM[851] = input_vector[106] << 4;
assign MEM[852] = input_vector[106] << 3;
assign MEM[853] = input_vector[106] << 2;
assign MEM[854] = input_vector[106] << 1;
assign MEM[855] = input_vector[106] << 0;
assign MEM[856] = -(input_vector[107] << 7);
assign MEM[857] = input_vector[107] << 6;
assign MEM[858] = input_vector[107] << 5;
assign MEM[859] = input_vector[107] << 4;
assign MEM[860] = input_vector[107] << 3;
assign MEM[861] = input_vector[107] << 2;
assign MEM[862] = input_vector[107] << 1;
assign MEM[863] = input_vector[107] << 0;
assign MEM[864] = -(input_vector[108] << 7);
assign MEM[865] = input_vector[108] << 6;
assign MEM[866] = input_vector[108] << 5;
assign MEM[867] = input_vector[108] << 4;
assign MEM[868] = input_vector[108] << 3;
assign MEM[869] = input_vector[108] << 2;
assign MEM[870] = input_vector[108] << 1;
assign MEM[871] = input_vector[108] << 0;
assign MEM[872] = -(input_vector[109] << 7);
assign MEM[873] = input_vector[109] << 6;
assign MEM[874] = input_vector[109] << 5;
assign MEM[875] = input_vector[109] << 4;
assign MEM[876] = input_vector[109] << 3;
assign MEM[877] = input_vector[109] << 2;
assign MEM[878] = input_vector[109] << 1;
assign MEM[879] = input_vector[109] << 0;
assign MEM[880] = -(input_vector[110] << 7);
assign MEM[881] = input_vector[110] << 6;
assign MEM[882] = input_vector[110] << 5;
assign MEM[883] = input_vector[110] << 4;
assign MEM[884] = input_vector[110] << 3;
assign MEM[885] = input_vector[110] << 2;
assign MEM[886] = input_vector[110] << 1;
assign MEM[887] = input_vector[110] << 0;
assign MEM[888] = -(input_vector[111] << 7);
assign MEM[889] = input_vector[111] << 6;
assign MEM[890] = input_vector[111] << 5;
assign MEM[891] = input_vector[111] << 4;
assign MEM[892] = input_vector[111] << 3;
assign MEM[893] = input_vector[111] << 2;
assign MEM[894] = input_vector[111] << 1;
assign MEM[895] = input_vector[111] << 0;
assign MEM[896] = -(input_vector[112] << 7);
assign MEM[897] = input_vector[112] << 6;
assign MEM[898] = input_vector[112] << 5;
assign MEM[899] = input_vector[112] << 4;
assign MEM[900] = input_vector[112] << 3;
assign MEM[901] = input_vector[112] << 2;
assign MEM[902] = input_vector[112] << 1;
assign MEM[903] = input_vector[112] << 0;
assign MEM[904] = -(input_vector[113] << 7);
assign MEM[905] = input_vector[113] << 6;
assign MEM[906] = input_vector[113] << 5;
assign MEM[907] = input_vector[113] << 4;
assign MEM[908] = input_vector[113] << 3;
assign MEM[909] = input_vector[113] << 2;
assign MEM[910] = input_vector[113] << 1;
assign MEM[911] = input_vector[113] << 0;
assign MEM[912] = -(input_vector[114] << 7);
assign MEM[913] = input_vector[114] << 6;
assign MEM[914] = input_vector[114] << 5;
assign MEM[915] = input_vector[114] << 4;
assign MEM[916] = input_vector[114] << 3;
assign MEM[917] = input_vector[114] << 2;
assign MEM[918] = input_vector[114] << 1;
assign MEM[919] = input_vector[114] << 0;
assign MEM[920] = -(input_vector[115] << 7);
assign MEM[921] = input_vector[115] << 6;
assign MEM[922] = input_vector[115] << 5;
assign MEM[923] = input_vector[115] << 4;
assign MEM[924] = input_vector[115] << 3;
assign MEM[925] = input_vector[115] << 2;
assign MEM[926] = input_vector[115] << 1;
assign MEM[927] = input_vector[115] << 0;
assign MEM[928] = -(input_vector[116] << 7);
assign MEM[929] = input_vector[116] << 6;
assign MEM[930] = input_vector[116] << 5;
assign MEM[931] = input_vector[116] << 4;
assign MEM[932] = input_vector[116] << 3;
assign MEM[933] = input_vector[116] << 2;
assign MEM[934] = input_vector[116] << 1;
assign MEM[935] = input_vector[116] << 0;
assign MEM[936] = -(input_vector[117] << 7);
assign MEM[937] = input_vector[117] << 6;
assign MEM[938] = input_vector[117] << 5;
assign MEM[939] = input_vector[117] << 4;
assign MEM[940] = input_vector[117] << 3;
assign MEM[941] = input_vector[117] << 2;
assign MEM[942] = input_vector[117] << 1;
assign MEM[943] = input_vector[117] << 0;
assign MEM[944] = -(input_vector[118] << 7);
assign MEM[945] = input_vector[118] << 6;
assign MEM[946] = input_vector[118] << 5;
assign MEM[947] = input_vector[118] << 4;
assign MEM[948] = input_vector[118] << 3;
assign MEM[949] = input_vector[118] << 2;
assign MEM[950] = input_vector[118] << 1;
assign MEM[951] = input_vector[118] << 0;
assign MEM[952] = -(input_vector[119] << 7);
assign MEM[953] = input_vector[119] << 6;
assign MEM[954] = input_vector[119] << 5;
assign MEM[955] = input_vector[119] << 4;
assign MEM[956] = input_vector[119] << 3;
assign MEM[957] = input_vector[119] << 2;
assign MEM[958] = input_vector[119] << 1;
assign MEM[959] = input_vector[119] << 0;
assign MEM[960] = -(input_vector[120] << 7);
assign MEM[961] = input_vector[120] << 6;
assign MEM[962] = input_vector[120] << 5;
assign MEM[963] = input_vector[120] << 4;
assign MEM[964] = input_vector[120] << 3;
assign MEM[965] = input_vector[120] << 2;
assign MEM[966] = input_vector[120] << 1;
assign MEM[967] = input_vector[120] << 0;
assign MEM[968] = -(input_vector[121] << 7);
assign MEM[969] = input_vector[121] << 6;
assign MEM[970] = input_vector[121] << 5;
assign MEM[971] = input_vector[121] << 4;
assign MEM[972] = input_vector[121] << 3;
assign MEM[973] = input_vector[121] << 2;
assign MEM[974] = input_vector[121] << 1;
assign MEM[975] = input_vector[121] << 0;
assign MEM[976] = -(input_vector[122] << 7);
assign MEM[977] = input_vector[122] << 6;
assign MEM[978] = input_vector[122] << 5;
assign MEM[979] = input_vector[122] << 4;
assign MEM[980] = input_vector[122] << 3;
assign MEM[981] = input_vector[122] << 2;
assign MEM[982] = input_vector[122] << 1;
assign MEM[983] = input_vector[122] << 0;
assign MEM[984] = -(input_vector[123] << 7);
assign MEM[985] = input_vector[123] << 6;
assign MEM[986] = input_vector[123] << 5;
assign MEM[987] = input_vector[123] << 4;
assign MEM[988] = input_vector[123] << 3;
assign MEM[989] = input_vector[123] << 2;
assign MEM[990] = input_vector[123] << 1;
assign MEM[991] = input_vector[123] << 0;
assign MEM[992] = -(input_vector[124] << 7);
assign MEM[993] = input_vector[124] << 6;
assign MEM[994] = input_vector[124] << 5;
assign MEM[995] = input_vector[124] << 4;
assign MEM[996] = input_vector[124] << 3;
assign MEM[997] = input_vector[124] << 2;
assign MEM[998] = input_vector[124] << 1;
assign MEM[999] = input_vector[124] << 0;
assign MEM[1000] = -(input_vector[125] << 7);
assign MEM[1001] = input_vector[125] << 6;
assign MEM[1002] = input_vector[125] << 5;
assign MEM[1003] = input_vector[125] << 4;
assign MEM[1004] = input_vector[125] << 3;
assign MEM[1005] = input_vector[125] << 2;
assign MEM[1006] = input_vector[125] << 1;
assign MEM[1007] = input_vector[125] << 0;
assign MEM[1008] = -(input_vector[126] << 7);
assign MEM[1009] = input_vector[126] << 6;
assign MEM[1010] = input_vector[126] << 5;
assign MEM[1011] = input_vector[126] << 4;
assign MEM[1012] = input_vector[126] << 3;
assign MEM[1013] = input_vector[126] << 2;
assign MEM[1014] = input_vector[126] << 1;
assign MEM[1015] = input_vector[126] << 0;
assign MEM[1016] = -(input_vector[127] << 7);
assign MEM[1017] = input_vector[127] << 6;
assign MEM[1018] = input_vector[127] << 5;
assign MEM[1019] = input_vector[127] << 4;
assign MEM[1020] = input_vector[127] << 3;
assign MEM[1021] = input_vector[127] << 2;
assign MEM[1022] = input_vector[127] << 1;
assign MEM[1023] = input_vector[127] << 0;
assign MEM[1024] = -(input_vector[128] << 7);
assign MEM[1025] = input_vector[128] << 6;
assign MEM[1026] = input_vector[128] << 5;
assign MEM[1027] = input_vector[128] << 4;
assign MEM[1028] = input_vector[128] << 3;
assign MEM[1029] = input_vector[128] << 2;
assign MEM[1030] = input_vector[128] << 1;
assign MEM[1031] = input_vector[128] << 0;
assign MEM[1032] = -(input_vector[129] << 7);
assign MEM[1033] = input_vector[129] << 6;
assign MEM[1034] = input_vector[129] << 5;
assign MEM[1035] = input_vector[129] << 4;
assign MEM[1036] = input_vector[129] << 3;
assign MEM[1037] = input_vector[129] << 2;
assign MEM[1038] = input_vector[129] << 1;
assign MEM[1039] = input_vector[129] << 0;
assign MEM[1040] = -(input_vector[130] << 7);
assign MEM[1041] = input_vector[130] << 6;
assign MEM[1042] = input_vector[130] << 5;
assign MEM[1043] = input_vector[130] << 4;
assign MEM[1044] = input_vector[130] << 3;
assign MEM[1045] = input_vector[130] << 2;
assign MEM[1046] = input_vector[130] << 1;
assign MEM[1047] = input_vector[130] << 0;
assign MEM[1048] = -(input_vector[131] << 7);
assign MEM[1049] = input_vector[131] << 6;
assign MEM[1050] = input_vector[131] << 5;
assign MEM[1051] = input_vector[131] << 4;
assign MEM[1052] = input_vector[131] << 3;
assign MEM[1053] = input_vector[131] << 2;
assign MEM[1054] = input_vector[131] << 1;
assign MEM[1055] = input_vector[131] << 0;
assign MEM[1056] = -(input_vector[132] << 7);
assign MEM[1057] = input_vector[132] << 6;
assign MEM[1058] = input_vector[132] << 5;
assign MEM[1059] = input_vector[132] << 4;
assign MEM[1060] = input_vector[132] << 3;
assign MEM[1061] = input_vector[132] << 2;
assign MEM[1062] = input_vector[132] << 1;
assign MEM[1063] = input_vector[132] << 0;
assign MEM[1064] = -(input_vector[133] << 7);
assign MEM[1065] = input_vector[133] << 6;
assign MEM[1066] = input_vector[133] << 5;
assign MEM[1067] = input_vector[133] << 4;
assign MEM[1068] = input_vector[133] << 3;
assign MEM[1069] = input_vector[133] << 2;
assign MEM[1070] = input_vector[133] << 1;
assign MEM[1071] = input_vector[133] << 0;
assign MEM[1072] = -(input_vector[134] << 7);
assign MEM[1073] = input_vector[134] << 6;
assign MEM[1074] = input_vector[134] << 5;
assign MEM[1075] = input_vector[134] << 4;
assign MEM[1076] = input_vector[134] << 3;
assign MEM[1077] = input_vector[134] << 2;
assign MEM[1078] = input_vector[134] << 1;
assign MEM[1079] = input_vector[134] << 0;
assign MEM[1080] = -(input_vector[135] << 7);
assign MEM[1081] = input_vector[135] << 6;
assign MEM[1082] = input_vector[135] << 5;
assign MEM[1083] = input_vector[135] << 4;
assign MEM[1084] = input_vector[135] << 3;
assign MEM[1085] = input_vector[135] << 2;
assign MEM[1086] = input_vector[135] << 1;
assign MEM[1087] = input_vector[135] << 0;
assign MEM[1088] = -(input_vector[136] << 7);
assign MEM[1089] = input_vector[136] << 6;
assign MEM[1090] = input_vector[136] << 5;
assign MEM[1091] = input_vector[136] << 4;
assign MEM[1092] = input_vector[136] << 3;
assign MEM[1093] = input_vector[136] << 2;
assign MEM[1094] = input_vector[136] << 1;
assign MEM[1095] = input_vector[136] << 0;
assign MEM[1096] = -(input_vector[137] << 7);
assign MEM[1097] = input_vector[137] << 6;
assign MEM[1098] = input_vector[137] << 5;
assign MEM[1099] = input_vector[137] << 4;
assign MEM[1100] = input_vector[137] << 3;
assign MEM[1101] = input_vector[137] << 2;
assign MEM[1102] = input_vector[137] << 1;
assign MEM[1103] = input_vector[137] << 0;
assign MEM[1104] = -(input_vector[138] << 7);
assign MEM[1105] = input_vector[138] << 6;
assign MEM[1106] = input_vector[138] << 5;
assign MEM[1107] = input_vector[138] << 4;
assign MEM[1108] = input_vector[138] << 3;
assign MEM[1109] = input_vector[138] << 2;
assign MEM[1110] = input_vector[138] << 1;
assign MEM[1111] = input_vector[138] << 0;
assign MEM[1112] = -(input_vector[139] << 7);
assign MEM[1113] = input_vector[139] << 6;
assign MEM[1114] = input_vector[139] << 5;
assign MEM[1115] = input_vector[139] << 4;
assign MEM[1116] = input_vector[139] << 3;
assign MEM[1117] = input_vector[139] << 2;
assign MEM[1118] = input_vector[139] << 1;
assign MEM[1119] = input_vector[139] << 0;
assign MEM[1120] = -(input_vector[140] << 7);
assign MEM[1121] = input_vector[140] << 6;
assign MEM[1122] = input_vector[140] << 5;
assign MEM[1123] = input_vector[140] << 4;
assign MEM[1124] = input_vector[140] << 3;
assign MEM[1125] = input_vector[140] << 2;
assign MEM[1126] = input_vector[140] << 1;
assign MEM[1127] = input_vector[140] << 0;
assign MEM[1128] = -(input_vector[141] << 7);
assign MEM[1129] = input_vector[141] << 6;
assign MEM[1130] = input_vector[141] << 5;
assign MEM[1131] = input_vector[141] << 4;
assign MEM[1132] = input_vector[141] << 3;
assign MEM[1133] = input_vector[141] << 2;
assign MEM[1134] = input_vector[141] << 1;
assign MEM[1135] = input_vector[141] << 0;
assign MEM[1136] = -(input_vector[142] << 7);
assign MEM[1137] = input_vector[142] << 6;
assign MEM[1138] = input_vector[142] << 5;
assign MEM[1139] = input_vector[142] << 4;
assign MEM[1140] = input_vector[142] << 3;
assign MEM[1141] = input_vector[142] << 2;
assign MEM[1142] = input_vector[142] << 1;
assign MEM[1143] = input_vector[142] << 0;
assign MEM[1144] = -(input_vector[143] << 7);
assign MEM[1145] = input_vector[143] << 6;
assign MEM[1146] = input_vector[143] << 5;
assign MEM[1147] = input_vector[143] << 4;
assign MEM[1148] = input_vector[143] << 3;
assign MEM[1149] = input_vector[143] << 2;
assign MEM[1150] = input_vector[143] << 1;
assign MEM[1151] = input_vector[143] << 0;
assign MEM[1152] = -(input_vector[144] << 7);
assign MEM[1153] = input_vector[144] << 6;
assign MEM[1154] = input_vector[144] << 5;
assign MEM[1155] = input_vector[144] << 4;
assign MEM[1156] = input_vector[144] << 3;
assign MEM[1157] = input_vector[144] << 2;
assign MEM[1158] = input_vector[144] << 1;
assign MEM[1159] = input_vector[144] << 0;
assign MEM[1160] = -(input_vector[145] << 7);
assign MEM[1161] = input_vector[145] << 6;
assign MEM[1162] = input_vector[145] << 5;
assign MEM[1163] = input_vector[145] << 4;
assign MEM[1164] = input_vector[145] << 3;
assign MEM[1165] = input_vector[145] << 2;
assign MEM[1166] = input_vector[145] << 1;
assign MEM[1167] = input_vector[145] << 0;
assign MEM[1168] = -(input_vector[146] << 7);
assign MEM[1169] = input_vector[146] << 6;
assign MEM[1170] = input_vector[146] << 5;
assign MEM[1171] = input_vector[146] << 4;
assign MEM[1172] = input_vector[146] << 3;
assign MEM[1173] = input_vector[146] << 2;
assign MEM[1174] = input_vector[146] << 1;
assign MEM[1175] = input_vector[146] << 0;
assign MEM[1176] = -(input_vector[147] << 7);
assign MEM[1177] = input_vector[147] << 6;
assign MEM[1178] = input_vector[147] << 5;
assign MEM[1179] = input_vector[147] << 4;
assign MEM[1180] = input_vector[147] << 3;
assign MEM[1181] = input_vector[147] << 2;
assign MEM[1182] = input_vector[147] << 1;
assign MEM[1183] = input_vector[147] << 0;
assign MEM[1184] = -(input_vector[148] << 7);
assign MEM[1185] = input_vector[148] << 6;
assign MEM[1186] = input_vector[148] << 5;
assign MEM[1187] = input_vector[148] << 4;
assign MEM[1188] = input_vector[148] << 3;
assign MEM[1189] = input_vector[148] << 2;
assign MEM[1190] = input_vector[148] << 1;
assign MEM[1191] = input_vector[148] << 0;
assign MEM[1192] = -(input_vector[149] << 7);
assign MEM[1193] = input_vector[149] << 6;
assign MEM[1194] = input_vector[149] << 5;
assign MEM[1195] = input_vector[149] << 4;
assign MEM[1196] = input_vector[149] << 3;
assign MEM[1197] = input_vector[149] << 2;
assign MEM[1198] = input_vector[149] << 1;
assign MEM[1199] = input_vector[149] << 0;
assign MEM[1200] = -(input_vector[150] << 7);
assign MEM[1201] = input_vector[150] << 6;
assign MEM[1202] = input_vector[150] << 5;
assign MEM[1203] = input_vector[150] << 4;
assign MEM[1204] = input_vector[150] << 3;
assign MEM[1205] = input_vector[150] << 2;
assign MEM[1206] = input_vector[150] << 1;
assign MEM[1207] = input_vector[150] << 0;
assign MEM[1208] = -(input_vector[151] << 7);
assign MEM[1209] = input_vector[151] << 6;
assign MEM[1210] = input_vector[151] << 5;
assign MEM[1211] = input_vector[151] << 4;
assign MEM[1212] = input_vector[151] << 3;
assign MEM[1213] = input_vector[151] << 2;
assign MEM[1214] = input_vector[151] << 1;
assign MEM[1215] = input_vector[151] << 0;
assign MEM[1216] = -(input_vector[152] << 7);
assign MEM[1217] = input_vector[152] << 6;
assign MEM[1218] = input_vector[152] << 5;
assign MEM[1219] = input_vector[152] << 4;
assign MEM[1220] = input_vector[152] << 3;
assign MEM[1221] = input_vector[152] << 2;
assign MEM[1222] = input_vector[152] << 1;
assign MEM[1223] = input_vector[152] << 0;
assign MEM[1224] = -(input_vector[153] << 7);
assign MEM[1225] = input_vector[153] << 6;
assign MEM[1226] = input_vector[153] << 5;
assign MEM[1227] = input_vector[153] << 4;
assign MEM[1228] = input_vector[153] << 3;
assign MEM[1229] = input_vector[153] << 2;
assign MEM[1230] = input_vector[153] << 1;
assign MEM[1231] = input_vector[153] << 0;
assign MEM[1232] = -(input_vector[154] << 7);
assign MEM[1233] = input_vector[154] << 6;
assign MEM[1234] = input_vector[154] << 5;
assign MEM[1235] = input_vector[154] << 4;
assign MEM[1236] = input_vector[154] << 3;
assign MEM[1237] = input_vector[154] << 2;
assign MEM[1238] = input_vector[154] << 1;
assign MEM[1239] = input_vector[154] << 0;
assign MEM[1240] = -(input_vector[155] << 7);
assign MEM[1241] = input_vector[155] << 6;
assign MEM[1242] = input_vector[155] << 5;
assign MEM[1243] = input_vector[155] << 4;
assign MEM[1244] = input_vector[155] << 3;
assign MEM[1245] = input_vector[155] << 2;
assign MEM[1246] = input_vector[155] << 1;
assign MEM[1247] = input_vector[155] << 0;
assign MEM[1248] = -(input_vector[156] << 7);
assign MEM[1249] = input_vector[156] << 6;
assign MEM[1250] = input_vector[156] << 5;
assign MEM[1251] = input_vector[156] << 4;
assign MEM[1252] = input_vector[156] << 3;
assign MEM[1253] = input_vector[156] << 2;
assign MEM[1254] = input_vector[156] << 1;
assign MEM[1255] = input_vector[156] << 0;
assign MEM[1256] = -(input_vector[157] << 7);
assign MEM[1257] = input_vector[157] << 6;
assign MEM[1258] = input_vector[157] << 5;
assign MEM[1259] = input_vector[157] << 4;
assign MEM[1260] = input_vector[157] << 3;
assign MEM[1261] = input_vector[157] << 2;
assign MEM[1262] = input_vector[157] << 1;
assign MEM[1263] = input_vector[157] << 0;
assign MEM[1264] = -(input_vector[158] << 7);
assign MEM[1265] = input_vector[158] << 6;
assign MEM[1266] = input_vector[158] << 5;
assign MEM[1267] = input_vector[158] << 4;
assign MEM[1268] = input_vector[158] << 3;
assign MEM[1269] = input_vector[158] << 2;
assign MEM[1270] = input_vector[158] << 1;
assign MEM[1271] = input_vector[158] << 0;
assign MEM[1272] = -(input_vector[159] << 7);
assign MEM[1273] = input_vector[159] << 6;
assign MEM[1274] = input_vector[159] << 5;
assign MEM[1275] = input_vector[159] << 4;
assign MEM[1276] = input_vector[159] << 3;
assign MEM[1277] = input_vector[159] << 2;
assign MEM[1278] = input_vector[159] << 1;
assign MEM[1279] = input_vector[159] << 0;
assign MEM[1280] = -(input_vector[160] << 7);
assign MEM[1281] = input_vector[160] << 6;
assign MEM[1282] = input_vector[160] << 5;
assign MEM[1283] = input_vector[160] << 4;
assign MEM[1284] = input_vector[160] << 3;
assign MEM[1285] = input_vector[160] << 2;
assign MEM[1286] = input_vector[160] << 1;
assign MEM[1287] = input_vector[160] << 0;
assign MEM[1288] = -(input_vector[161] << 7);
assign MEM[1289] = input_vector[161] << 6;
assign MEM[1290] = input_vector[161] << 5;
assign MEM[1291] = input_vector[161] << 4;
assign MEM[1292] = input_vector[161] << 3;
assign MEM[1293] = input_vector[161] << 2;
assign MEM[1294] = input_vector[161] << 1;
assign MEM[1295] = input_vector[161] << 0;
assign MEM[1296] = -(input_vector[162] << 7);
assign MEM[1297] = input_vector[162] << 6;
assign MEM[1298] = input_vector[162] << 5;
assign MEM[1299] = input_vector[162] << 4;
assign MEM[1300] = input_vector[162] << 3;
assign MEM[1301] = input_vector[162] << 2;
assign MEM[1302] = input_vector[162] << 1;
assign MEM[1303] = input_vector[162] << 0;
assign MEM[1304] = -(input_vector[163] << 7);
assign MEM[1305] = input_vector[163] << 6;
assign MEM[1306] = input_vector[163] << 5;
assign MEM[1307] = input_vector[163] << 4;
assign MEM[1308] = input_vector[163] << 3;
assign MEM[1309] = input_vector[163] << 2;
assign MEM[1310] = input_vector[163] << 1;
assign MEM[1311] = input_vector[163] << 0;
assign MEM[1312] = -(input_vector[164] << 7);
assign MEM[1313] = input_vector[164] << 6;
assign MEM[1314] = input_vector[164] << 5;
assign MEM[1315] = input_vector[164] << 4;
assign MEM[1316] = input_vector[164] << 3;
assign MEM[1317] = input_vector[164] << 2;
assign MEM[1318] = input_vector[164] << 1;
assign MEM[1319] = input_vector[164] << 0;
assign MEM[1320] = -(input_vector[165] << 7);
assign MEM[1321] = input_vector[165] << 6;
assign MEM[1322] = input_vector[165] << 5;
assign MEM[1323] = input_vector[165] << 4;
assign MEM[1324] = input_vector[165] << 3;
assign MEM[1325] = input_vector[165] << 2;
assign MEM[1326] = input_vector[165] << 1;
assign MEM[1327] = input_vector[165] << 0;
assign MEM[1328] = -(input_vector[166] << 7);
assign MEM[1329] = input_vector[166] << 6;
assign MEM[1330] = input_vector[166] << 5;
assign MEM[1331] = input_vector[166] << 4;
assign MEM[1332] = input_vector[166] << 3;
assign MEM[1333] = input_vector[166] << 2;
assign MEM[1334] = input_vector[166] << 1;
assign MEM[1335] = input_vector[166] << 0;
assign MEM[1336] = -(input_vector[167] << 7);
assign MEM[1337] = input_vector[167] << 6;
assign MEM[1338] = input_vector[167] << 5;
assign MEM[1339] = input_vector[167] << 4;
assign MEM[1340] = input_vector[167] << 3;
assign MEM[1341] = input_vector[167] << 2;
assign MEM[1342] = input_vector[167] << 1;
assign MEM[1343] = input_vector[167] << 0;
assign MEM[1344] = -(input_vector[168] << 7);
assign MEM[1345] = input_vector[168] << 6;
assign MEM[1346] = input_vector[168] << 5;
assign MEM[1347] = input_vector[168] << 4;
assign MEM[1348] = input_vector[168] << 3;
assign MEM[1349] = input_vector[168] << 2;
assign MEM[1350] = input_vector[168] << 1;
assign MEM[1351] = input_vector[168] << 0;
assign MEM[1352] = -(input_vector[169] << 7);
assign MEM[1353] = input_vector[169] << 6;
assign MEM[1354] = input_vector[169] << 5;
assign MEM[1355] = input_vector[169] << 4;
assign MEM[1356] = input_vector[169] << 3;
assign MEM[1357] = input_vector[169] << 2;
assign MEM[1358] = input_vector[169] << 1;
assign MEM[1359] = input_vector[169] << 0;
assign MEM[1360] = -(input_vector[170] << 7);
assign MEM[1361] = input_vector[170] << 6;
assign MEM[1362] = input_vector[170] << 5;
assign MEM[1363] = input_vector[170] << 4;
assign MEM[1364] = input_vector[170] << 3;
assign MEM[1365] = input_vector[170] << 2;
assign MEM[1366] = input_vector[170] << 1;
assign MEM[1367] = input_vector[170] << 0;
assign MEM[1368] = -(input_vector[171] << 7);
assign MEM[1369] = input_vector[171] << 6;
assign MEM[1370] = input_vector[171] << 5;
assign MEM[1371] = input_vector[171] << 4;
assign MEM[1372] = input_vector[171] << 3;
assign MEM[1373] = input_vector[171] << 2;
assign MEM[1374] = input_vector[171] << 1;
assign MEM[1375] = input_vector[171] << 0;
assign MEM[1376] = -(input_vector[172] << 7);
assign MEM[1377] = input_vector[172] << 6;
assign MEM[1378] = input_vector[172] << 5;
assign MEM[1379] = input_vector[172] << 4;
assign MEM[1380] = input_vector[172] << 3;
assign MEM[1381] = input_vector[172] << 2;
assign MEM[1382] = input_vector[172] << 1;
assign MEM[1383] = input_vector[172] << 0;
assign MEM[1384] = -(input_vector[173] << 7);
assign MEM[1385] = input_vector[173] << 6;
assign MEM[1386] = input_vector[173] << 5;
assign MEM[1387] = input_vector[173] << 4;
assign MEM[1388] = input_vector[173] << 3;
assign MEM[1389] = input_vector[173] << 2;
assign MEM[1390] = input_vector[173] << 1;
assign MEM[1391] = input_vector[173] << 0;
assign MEM[1392] = -(input_vector[174] << 7);
assign MEM[1393] = input_vector[174] << 6;
assign MEM[1394] = input_vector[174] << 5;
assign MEM[1395] = input_vector[174] << 4;
assign MEM[1396] = input_vector[174] << 3;
assign MEM[1397] = input_vector[174] << 2;
assign MEM[1398] = input_vector[174] << 1;
assign MEM[1399] = input_vector[174] << 0;
assign MEM[1400] = -(input_vector[175] << 7);
assign MEM[1401] = input_vector[175] << 6;
assign MEM[1402] = input_vector[175] << 5;
assign MEM[1403] = input_vector[175] << 4;
assign MEM[1404] = input_vector[175] << 3;
assign MEM[1405] = input_vector[175] << 2;
assign MEM[1406] = input_vector[175] << 1;
assign MEM[1407] = input_vector[175] << 0;
assign MEM[1408] = -(input_vector[176] << 7);
assign MEM[1409] = input_vector[176] << 6;
assign MEM[1410] = input_vector[176] << 5;
assign MEM[1411] = input_vector[176] << 4;
assign MEM[1412] = input_vector[176] << 3;
assign MEM[1413] = input_vector[176] << 2;
assign MEM[1414] = input_vector[176] << 1;
assign MEM[1415] = input_vector[176] << 0;
assign MEM[1416] = -(input_vector[177] << 7);
assign MEM[1417] = input_vector[177] << 6;
assign MEM[1418] = input_vector[177] << 5;
assign MEM[1419] = input_vector[177] << 4;
assign MEM[1420] = input_vector[177] << 3;
assign MEM[1421] = input_vector[177] << 2;
assign MEM[1422] = input_vector[177] << 1;
assign MEM[1423] = input_vector[177] << 0;
assign MEM[1424] = -(input_vector[178] << 7);
assign MEM[1425] = input_vector[178] << 6;
assign MEM[1426] = input_vector[178] << 5;
assign MEM[1427] = input_vector[178] << 4;
assign MEM[1428] = input_vector[178] << 3;
assign MEM[1429] = input_vector[178] << 2;
assign MEM[1430] = input_vector[178] << 1;
assign MEM[1431] = input_vector[178] << 0;
assign MEM[1432] = -(input_vector[179] << 7);
assign MEM[1433] = input_vector[179] << 6;
assign MEM[1434] = input_vector[179] << 5;
assign MEM[1435] = input_vector[179] << 4;
assign MEM[1436] = input_vector[179] << 3;
assign MEM[1437] = input_vector[179] << 2;
assign MEM[1438] = input_vector[179] << 1;
assign MEM[1439] = input_vector[179] << 0;
assign MEM[1440] = -(input_vector[180] << 7);
assign MEM[1441] = input_vector[180] << 6;
assign MEM[1442] = input_vector[180] << 5;
assign MEM[1443] = input_vector[180] << 4;
assign MEM[1444] = input_vector[180] << 3;
assign MEM[1445] = input_vector[180] << 2;
assign MEM[1446] = input_vector[180] << 1;
assign MEM[1447] = input_vector[180] << 0;
assign MEM[1448] = -(input_vector[181] << 7);
assign MEM[1449] = input_vector[181] << 6;
assign MEM[1450] = input_vector[181] << 5;
assign MEM[1451] = input_vector[181] << 4;
assign MEM[1452] = input_vector[181] << 3;
assign MEM[1453] = input_vector[181] << 2;
assign MEM[1454] = input_vector[181] << 1;
assign MEM[1455] = input_vector[181] << 0;
assign MEM[1456] = -(input_vector[182] << 7);
assign MEM[1457] = input_vector[182] << 6;
assign MEM[1458] = input_vector[182] << 5;
assign MEM[1459] = input_vector[182] << 4;
assign MEM[1460] = input_vector[182] << 3;
assign MEM[1461] = input_vector[182] << 2;
assign MEM[1462] = input_vector[182] << 1;
assign MEM[1463] = input_vector[182] << 0;
assign MEM[1464] = -(input_vector[183] << 7);
assign MEM[1465] = input_vector[183] << 6;
assign MEM[1466] = input_vector[183] << 5;
assign MEM[1467] = input_vector[183] << 4;
assign MEM[1468] = input_vector[183] << 3;
assign MEM[1469] = input_vector[183] << 2;
assign MEM[1470] = input_vector[183] << 1;
assign MEM[1471] = input_vector[183] << 0;
assign MEM[1472] = -(input_vector[184] << 7);
assign MEM[1473] = input_vector[184] << 6;
assign MEM[1474] = input_vector[184] << 5;
assign MEM[1475] = input_vector[184] << 4;
assign MEM[1476] = input_vector[184] << 3;
assign MEM[1477] = input_vector[184] << 2;
assign MEM[1478] = input_vector[184] << 1;
assign MEM[1479] = input_vector[184] << 0;
assign MEM[1480] = -(input_vector[185] << 7);
assign MEM[1481] = input_vector[185] << 6;
assign MEM[1482] = input_vector[185] << 5;
assign MEM[1483] = input_vector[185] << 4;
assign MEM[1484] = input_vector[185] << 3;
assign MEM[1485] = input_vector[185] << 2;
assign MEM[1486] = input_vector[185] << 1;
assign MEM[1487] = input_vector[185] << 0;
assign MEM[1488] = -(input_vector[186] << 7);
assign MEM[1489] = input_vector[186] << 6;
assign MEM[1490] = input_vector[186] << 5;
assign MEM[1491] = input_vector[186] << 4;
assign MEM[1492] = input_vector[186] << 3;
assign MEM[1493] = input_vector[186] << 2;
assign MEM[1494] = input_vector[186] << 1;
assign MEM[1495] = input_vector[186] << 0;
assign MEM[1496] = -(input_vector[187] << 7);
assign MEM[1497] = input_vector[187] << 6;
assign MEM[1498] = input_vector[187] << 5;
assign MEM[1499] = input_vector[187] << 4;
assign MEM[1500] = input_vector[187] << 3;
assign MEM[1501] = input_vector[187] << 2;
assign MEM[1502] = input_vector[187] << 1;
assign MEM[1503] = input_vector[187] << 0;
assign MEM[1504] = -(input_vector[188] << 7);
assign MEM[1505] = input_vector[188] << 6;
assign MEM[1506] = input_vector[188] << 5;
assign MEM[1507] = input_vector[188] << 4;
assign MEM[1508] = input_vector[188] << 3;
assign MEM[1509] = input_vector[188] << 2;
assign MEM[1510] = input_vector[188] << 1;
assign MEM[1511] = input_vector[188] << 0;
assign MEM[1512] = -(input_vector[189] << 7);
assign MEM[1513] = input_vector[189] << 6;
assign MEM[1514] = input_vector[189] << 5;
assign MEM[1515] = input_vector[189] << 4;
assign MEM[1516] = input_vector[189] << 3;
assign MEM[1517] = input_vector[189] << 2;
assign MEM[1518] = input_vector[189] << 1;
assign MEM[1519] = input_vector[189] << 0;
assign MEM[1520] = -(input_vector[190] << 7);
assign MEM[1521] = input_vector[190] << 6;
assign MEM[1522] = input_vector[190] << 5;
assign MEM[1523] = input_vector[190] << 4;
assign MEM[1524] = input_vector[190] << 3;
assign MEM[1525] = input_vector[190] << 2;
assign MEM[1526] = input_vector[190] << 1;
assign MEM[1527] = input_vector[190] << 0;
assign MEM[1528] = -(input_vector[191] << 7);
assign MEM[1529] = input_vector[191] << 6;
assign MEM[1530] = input_vector[191] << 5;
assign MEM[1531] = input_vector[191] << 4;
assign MEM[1532] = input_vector[191] << 3;
assign MEM[1533] = input_vector[191] << 2;
assign MEM[1534] = input_vector[191] << 1;
assign MEM[1535] = input_vector[191] << 0;
assign MEM[1536] = -(input_vector[192] << 7);
assign MEM[1537] = input_vector[192] << 6;
assign MEM[1538] = input_vector[192] << 5;
assign MEM[1539] = input_vector[192] << 4;
assign MEM[1540] = input_vector[192] << 3;
assign MEM[1541] = input_vector[192] << 2;
assign MEM[1542] = input_vector[192] << 1;
assign MEM[1543] = input_vector[192] << 0;
assign MEM[1544] = -(input_vector[193] << 7);
assign MEM[1545] = input_vector[193] << 6;
assign MEM[1546] = input_vector[193] << 5;
assign MEM[1547] = input_vector[193] << 4;
assign MEM[1548] = input_vector[193] << 3;
assign MEM[1549] = input_vector[193] << 2;
assign MEM[1550] = input_vector[193] << 1;
assign MEM[1551] = input_vector[193] << 0;
assign MEM[1552] = -(input_vector[194] << 7);
assign MEM[1553] = input_vector[194] << 6;
assign MEM[1554] = input_vector[194] << 5;
assign MEM[1555] = input_vector[194] << 4;
assign MEM[1556] = input_vector[194] << 3;
assign MEM[1557] = input_vector[194] << 2;
assign MEM[1558] = input_vector[194] << 1;
assign MEM[1559] = input_vector[194] << 0;
assign MEM[1560] = -(input_vector[195] << 7);
assign MEM[1561] = input_vector[195] << 6;
assign MEM[1562] = input_vector[195] << 5;
assign MEM[1563] = input_vector[195] << 4;
assign MEM[1564] = input_vector[195] << 3;
assign MEM[1565] = input_vector[195] << 2;
assign MEM[1566] = input_vector[195] << 1;
assign MEM[1567] = input_vector[195] << 0;
assign MEM[1568] = -(input_vector[196] << 7);
assign MEM[1569] = input_vector[196] << 6;
assign MEM[1570] = input_vector[196] << 5;
assign MEM[1571] = input_vector[196] << 4;
assign MEM[1572] = input_vector[196] << 3;
assign MEM[1573] = input_vector[196] << 2;
assign MEM[1574] = input_vector[196] << 1;
assign MEM[1575] = input_vector[196] << 0;
assign MEM[1576] = -(input_vector[197] << 7);
assign MEM[1577] = input_vector[197] << 6;
assign MEM[1578] = input_vector[197] << 5;
assign MEM[1579] = input_vector[197] << 4;
assign MEM[1580] = input_vector[197] << 3;
assign MEM[1581] = input_vector[197] << 2;
assign MEM[1582] = input_vector[197] << 1;
assign MEM[1583] = input_vector[197] << 0;
assign MEM[1584] = -(input_vector[198] << 7);
assign MEM[1585] = input_vector[198] << 6;
assign MEM[1586] = input_vector[198] << 5;
assign MEM[1587] = input_vector[198] << 4;
assign MEM[1588] = input_vector[198] << 3;
assign MEM[1589] = input_vector[198] << 2;
assign MEM[1590] = input_vector[198] << 1;
assign MEM[1591] = input_vector[198] << 0;
assign MEM[1592] = -(input_vector[199] << 7);
assign MEM[1593] = input_vector[199] << 6;
assign MEM[1594] = input_vector[199] << 5;
assign MEM[1595] = input_vector[199] << 4;
assign MEM[1596] = input_vector[199] << 3;
assign MEM[1597] = input_vector[199] << 2;
assign MEM[1598] = input_vector[199] << 1;
assign MEM[1599] = input_vector[199] << 0;
assign MEM[1600] = -(input_vector[200] << 7);
assign MEM[1601] = input_vector[200] << 6;
assign MEM[1602] = input_vector[200] << 5;
assign MEM[1603] = input_vector[200] << 4;
assign MEM[1604] = input_vector[200] << 3;
assign MEM[1605] = input_vector[200] << 2;
assign MEM[1606] = input_vector[200] << 1;
assign MEM[1607] = input_vector[200] << 0;
assign MEM[1608] = -(input_vector[201] << 7);
assign MEM[1609] = input_vector[201] << 6;
assign MEM[1610] = input_vector[201] << 5;
assign MEM[1611] = input_vector[201] << 4;
assign MEM[1612] = input_vector[201] << 3;
assign MEM[1613] = input_vector[201] << 2;
assign MEM[1614] = input_vector[201] << 1;
assign MEM[1615] = input_vector[201] << 0;
assign MEM[1616] = -(input_vector[202] << 7);
assign MEM[1617] = input_vector[202] << 6;
assign MEM[1618] = input_vector[202] << 5;
assign MEM[1619] = input_vector[202] << 4;
assign MEM[1620] = input_vector[202] << 3;
assign MEM[1621] = input_vector[202] << 2;
assign MEM[1622] = input_vector[202] << 1;
assign MEM[1623] = input_vector[202] << 0;
assign MEM[1624] = -(input_vector[203] << 7);
assign MEM[1625] = input_vector[203] << 6;
assign MEM[1626] = input_vector[203] << 5;
assign MEM[1627] = input_vector[203] << 4;
assign MEM[1628] = input_vector[203] << 3;
assign MEM[1629] = input_vector[203] << 2;
assign MEM[1630] = input_vector[203] << 1;
assign MEM[1631] = input_vector[203] << 0;
assign MEM[1632] = -(input_vector[204] << 7);
assign MEM[1633] = input_vector[204] << 6;
assign MEM[1634] = input_vector[204] << 5;
assign MEM[1635] = input_vector[204] << 4;
assign MEM[1636] = input_vector[204] << 3;
assign MEM[1637] = input_vector[204] << 2;
assign MEM[1638] = input_vector[204] << 1;
assign MEM[1639] = input_vector[204] << 0;
assign MEM[1640] = -(input_vector[205] << 7);
assign MEM[1641] = input_vector[205] << 6;
assign MEM[1642] = input_vector[205] << 5;
assign MEM[1643] = input_vector[205] << 4;
assign MEM[1644] = input_vector[205] << 3;
assign MEM[1645] = input_vector[205] << 2;
assign MEM[1646] = input_vector[205] << 1;
assign MEM[1647] = input_vector[205] << 0;
assign MEM[1648] = -(input_vector[206] << 7);
assign MEM[1649] = input_vector[206] << 6;
assign MEM[1650] = input_vector[206] << 5;
assign MEM[1651] = input_vector[206] << 4;
assign MEM[1652] = input_vector[206] << 3;
assign MEM[1653] = input_vector[206] << 2;
assign MEM[1654] = input_vector[206] << 1;
assign MEM[1655] = input_vector[206] << 0;
assign MEM[1656] = -(input_vector[207] << 7);
assign MEM[1657] = input_vector[207] << 6;
assign MEM[1658] = input_vector[207] << 5;
assign MEM[1659] = input_vector[207] << 4;
assign MEM[1660] = input_vector[207] << 3;
assign MEM[1661] = input_vector[207] << 2;
assign MEM[1662] = input_vector[207] << 1;
assign MEM[1663] = input_vector[207] << 0;
assign MEM[1664] = -(input_vector[208] << 7);
assign MEM[1665] = input_vector[208] << 6;
assign MEM[1666] = input_vector[208] << 5;
assign MEM[1667] = input_vector[208] << 4;
assign MEM[1668] = input_vector[208] << 3;
assign MEM[1669] = input_vector[208] << 2;
assign MEM[1670] = input_vector[208] << 1;
assign MEM[1671] = input_vector[208] << 0;
assign MEM[1672] = -(input_vector[209] << 7);
assign MEM[1673] = input_vector[209] << 6;
assign MEM[1674] = input_vector[209] << 5;
assign MEM[1675] = input_vector[209] << 4;
assign MEM[1676] = input_vector[209] << 3;
assign MEM[1677] = input_vector[209] << 2;
assign MEM[1678] = input_vector[209] << 1;
assign MEM[1679] = input_vector[209] << 0;
assign MEM[1680] = -(input_vector[210] << 7);
assign MEM[1681] = input_vector[210] << 6;
assign MEM[1682] = input_vector[210] << 5;
assign MEM[1683] = input_vector[210] << 4;
assign MEM[1684] = input_vector[210] << 3;
assign MEM[1685] = input_vector[210] << 2;
assign MEM[1686] = input_vector[210] << 1;
assign MEM[1687] = input_vector[210] << 0;
assign MEM[1688] = -(input_vector[211] << 7);
assign MEM[1689] = input_vector[211] << 6;
assign MEM[1690] = input_vector[211] << 5;
assign MEM[1691] = input_vector[211] << 4;
assign MEM[1692] = input_vector[211] << 3;
assign MEM[1693] = input_vector[211] << 2;
assign MEM[1694] = input_vector[211] << 1;
assign MEM[1695] = input_vector[211] << 0;
assign MEM[1696] = -(input_vector[212] << 7);
assign MEM[1697] = input_vector[212] << 6;
assign MEM[1698] = input_vector[212] << 5;
assign MEM[1699] = input_vector[212] << 4;
assign MEM[1700] = input_vector[212] << 3;
assign MEM[1701] = input_vector[212] << 2;
assign MEM[1702] = input_vector[212] << 1;
assign MEM[1703] = input_vector[212] << 0;
assign MEM[1704] = -(input_vector[213] << 7);
assign MEM[1705] = input_vector[213] << 6;
assign MEM[1706] = input_vector[213] << 5;
assign MEM[1707] = input_vector[213] << 4;
assign MEM[1708] = input_vector[213] << 3;
assign MEM[1709] = input_vector[213] << 2;
assign MEM[1710] = input_vector[213] << 1;
assign MEM[1711] = input_vector[213] << 0;
assign MEM[1712] = -(input_vector[214] << 7);
assign MEM[1713] = input_vector[214] << 6;
assign MEM[1714] = input_vector[214] << 5;
assign MEM[1715] = input_vector[214] << 4;
assign MEM[1716] = input_vector[214] << 3;
assign MEM[1717] = input_vector[214] << 2;
assign MEM[1718] = input_vector[214] << 1;
assign MEM[1719] = input_vector[214] << 0;
assign MEM[1720] = -(input_vector[215] << 7);
assign MEM[1721] = input_vector[215] << 6;
assign MEM[1722] = input_vector[215] << 5;
assign MEM[1723] = input_vector[215] << 4;
assign MEM[1724] = input_vector[215] << 3;
assign MEM[1725] = input_vector[215] << 2;
assign MEM[1726] = input_vector[215] << 1;
assign MEM[1727] = input_vector[215] << 0;
assign MEM[1728] = -(input_vector[216] << 7);
assign MEM[1729] = input_vector[216] << 6;
assign MEM[1730] = input_vector[216] << 5;
assign MEM[1731] = input_vector[216] << 4;
assign MEM[1732] = input_vector[216] << 3;
assign MEM[1733] = input_vector[216] << 2;
assign MEM[1734] = input_vector[216] << 1;
assign MEM[1735] = input_vector[216] << 0;
assign MEM[1736] = -(input_vector[217] << 7);
assign MEM[1737] = input_vector[217] << 6;
assign MEM[1738] = input_vector[217] << 5;
assign MEM[1739] = input_vector[217] << 4;
assign MEM[1740] = input_vector[217] << 3;
assign MEM[1741] = input_vector[217] << 2;
assign MEM[1742] = input_vector[217] << 1;
assign MEM[1743] = input_vector[217] << 0;
assign MEM[1744] = -(input_vector[218] << 7);
assign MEM[1745] = input_vector[218] << 6;
assign MEM[1746] = input_vector[218] << 5;
assign MEM[1747] = input_vector[218] << 4;
assign MEM[1748] = input_vector[218] << 3;
assign MEM[1749] = input_vector[218] << 2;
assign MEM[1750] = input_vector[218] << 1;
assign MEM[1751] = input_vector[218] << 0;
assign MEM[1752] = -(input_vector[219] << 7);
assign MEM[1753] = input_vector[219] << 6;
assign MEM[1754] = input_vector[219] << 5;
assign MEM[1755] = input_vector[219] << 4;
assign MEM[1756] = input_vector[219] << 3;
assign MEM[1757] = input_vector[219] << 2;
assign MEM[1758] = input_vector[219] << 1;
assign MEM[1759] = input_vector[219] << 0;
assign MEM[1760] = -(input_vector[220] << 7);
assign MEM[1761] = input_vector[220] << 6;
assign MEM[1762] = input_vector[220] << 5;
assign MEM[1763] = input_vector[220] << 4;
assign MEM[1764] = input_vector[220] << 3;
assign MEM[1765] = input_vector[220] << 2;
assign MEM[1766] = input_vector[220] << 1;
assign MEM[1767] = input_vector[220] << 0;
assign MEM[1768] = -(input_vector[221] << 7);
assign MEM[1769] = input_vector[221] << 6;
assign MEM[1770] = input_vector[221] << 5;
assign MEM[1771] = input_vector[221] << 4;
assign MEM[1772] = input_vector[221] << 3;
assign MEM[1773] = input_vector[221] << 2;
assign MEM[1774] = input_vector[221] << 1;
assign MEM[1775] = input_vector[221] << 0;
assign MEM[1776] = -(input_vector[222] << 7);
assign MEM[1777] = input_vector[222] << 6;
assign MEM[1778] = input_vector[222] << 5;
assign MEM[1779] = input_vector[222] << 4;
assign MEM[1780] = input_vector[222] << 3;
assign MEM[1781] = input_vector[222] << 2;
assign MEM[1782] = input_vector[222] << 1;
assign MEM[1783] = input_vector[222] << 0;
assign MEM[1784] = -(input_vector[223] << 7);
assign MEM[1785] = input_vector[223] << 6;
assign MEM[1786] = input_vector[223] << 5;
assign MEM[1787] = input_vector[223] << 4;
assign MEM[1788] = input_vector[223] << 3;
assign MEM[1789] = input_vector[223] << 2;
assign MEM[1790] = input_vector[223] << 1;
assign MEM[1791] = input_vector[223] << 0;
assign MEM[1792] = -(input_vector[224] << 7);
assign MEM[1793] = input_vector[224] << 6;
assign MEM[1794] = input_vector[224] << 5;
assign MEM[1795] = input_vector[224] << 4;
assign MEM[1796] = input_vector[224] << 3;
assign MEM[1797] = input_vector[224] << 2;
assign MEM[1798] = input_vector[224] << 1;
assign MEM[1799] = input_vector[224] << 0;
assign MEM[1800] = -(input_vector[225] << 7);
assign MEM[1801] = input_vector[225] << 6;
assign MEM[1802] = input_vector[225] << 5;
assign MEM[1803] = input_vector[225] << 4;
assign MEM[1804] = input_vector[225] << 3;
assign MEM[1805] = input_vector[225] << 2;
assign MEM[1806] = input_vector[225] << 1;
assign MEM[1807] = input_vector[225] << 0;
assign MEM[1808] = -(input_vector[226] << 7);
assign MEM[1809] = input_vector[226] << 6;
assign MEM[1810] = input_vector[226] << 5;
assign MEM[1811] = input_vector[226] << 4;
assign MEM[1812] = input_vector[226] << 3;
assign MEM[1813] = input_vector[226] << 2;
assign MEM[1814] = input_vector[226] << 1;
assign MEM[1815] = input_vector[226] << 0;
assign MEM[1816] = -(input_vector[227] << 7);
assign MEM[1817] = input_vector[227] << 6;
assign MEM[1818] = input_vector[227] << 5;
assign MEM[1819] = input_vector[227] << 4;
assign MEM[1820] = input_vector[227] << 3;
assign MEM[1821] = input_vector[227] << 2;
assign MEM[1822] = input_vector[227] << 1;
assign MEM[1823] = input_vector[227] << 0;
assign MEM[1824] = -(input_vector[228] << 7);
assign MEM[1825] = input_vector[228] << 6;
assign MEM[1826] = input_vector[228] << 5;
assign MEM[1827] = input_vector[228] << 4;
assign MEM[1828] = input_vector[228] << 3;
assign MEM[1829] = input_vector[228] << 2;
assign MEM[1830] = input_vector[228] << 1;
assign MEM[1831] = input_vector[228] << 0;
assign MEM[1832] = -(input_vector[229] << 7);
assign MEM[1833] = input_vector[229] << 6;
assign MEM[1834] = input_vector[229] << 5;
assign MEM[1835] = input_vector[229] << 4;
assign MEM[1836] = input_vector[229] << 3;
assign MEM[1837] = input_vector[229] << 2;
assign MEM[1838] = input_vector[229] << 1;
assign MEM[1839] = input_vector[229] << 0;
assign MEM[1840] = -(input_vector[230] << 7);
assign MEM[1841] = input_vector[230] << 6;
assign MEM[1842] = input_vector[230] << 5;
assign MEM[1843] = input_vector[230] << 4;
assign MEM[1844] = input_vector[230] << 3;
assign MEM[1845] = input_vector[230] << 2;
assign MEM[1846] = input_vector[230] << 1;
assign MEM[1847] = input_vector[230] << 0;
assign MEM[1848] = -(input_vector[231] << 7);
assign MEM[1849] = input_vector[231] << 6;
assign MEM[1850] = input_vector[231] << 5;
assign MEM[1851] = input_vector[231] << 4;
assign MEM[1852] = input_vector[231] << 3;
assign MEM[1853] = input_vector[231] << 2;
assign MEM[1854] = input_vector[231] << 1;
assign MEM[1855] = input_vector[231] << 0;
assign MEM[1856] = -(input_vector[232] << 7);
assign MEM[1857] = input_vector[232] << 6;
assign MEM[1858] = input_vector[232] << 5;
assign MEM[1859] = input_vector[232] << 4;
assign MEM[1860] = input_vector[232] << 3;
assign MEM[1861] = input_vector[232] << 2;
assign MEM[1862] = input_vector[232] << 1;
assign MEM[1863] = input_vector[232] << 0;
assign MEM[1864] = -(input_vector[233] << 7);
assign MEM[1865] = input_vector[233] << 6;
assign MEM[1866] = input_vector[233] << 5;
assign MEM[1867] = input_vector[233] << 4;
assign MEM[1868] = input_vector[233] << 3;
assign MEM[1869] = input_vector[233] << 2;
assign MEM[1870] = input_vector[233] << 1;
assign MEM[1871] = input_vector[233] << 0;
assign MEM[1872] = -(input_vector[234] << 7);
assign MEM[1873] = input_vector[234] << 6;
assign MEM[1874] = input_vector[234] << 5;
assign MEM[1875] = input_vector[234] << 4;
assign MEM[1876] = input_vector[234] << 3;
assign MEM[1877] = input_vector[234] << 2;
assign MEM[1878] = input_vector[234] << 1;
assign MEM[1879] = input_vector[234] << 0;
assign MEM[1880] = -(input_vector[235] << 7);
assign MEM[1881] = input_vector[235] << 6;
assign MEM[1882] = input_vector[235] << 5;
assign MEM[1883] = input_vector[235] << 4;
assign MEM[1884] = input_vector[235] << 3;
assign MEM[1885] = input_vector[235] << 2;
assign MEM[1886] = input_vector[235] << 1;
assign MEM[1887] = input_vector[235] << 0;
assign MEM[1888] = -(input_vector[236] << 7);
assign MEM[1889] = input_vector[236] << 6;
assign MEM[1890] = input_vector[236] << 5;
assign MEM[1891] = input_vector[236] << 4;
assign MEM[1892] = input_vector[236] << 3;
assign MEM[1893] = input_vector[236] << 2;
assign MEM[1894] = input_vector[236] << 1;
assign MEM[1895] = input_vector[236] << 0;
assign MEM[1896] = -(input_vector[237] << 7);
assign MEM[1897] = input_vector[237] << 6;
assign MEM[1898] = input_vector[237] << 5;
assign MEM[1899] = input_vector[237] << 4;
assign MEM[1900] = input_vector[237] << 3;
assign MEM[1901] = input_vector[237] << 2;
assign MEM[1902] = input_vector[237] << 1;
assign MEM[1903] = input_vector[237] << 0;
assign MEM[1904] = -(input_vector[238] << 7);
assign MEM[1905] = input_vector[238] << 6;
assign MEM[1906] = input_vector[238] << 5;
assign MEM[1907] = input_vector[238] << 4;
assign MEM[1908] = input_vector[238] << 3;
assign MEM[1909] = input_vector[238] << 2;
assign MEM[1910] = input_vector[238] << 1;
assign MEM[1911] = input_vector[238] << 0;
assign MEM[1912] = -(input_vector[239] << 7);
assign MEM[1913] = input_vector[239] << 6;
assign MEM[1914] = input_vector[239] << 5;
assign MEM[1915] = input_vector[239] << 4;
assign MEM[1916] = input_vector[239] << 3;
assign MEM[1917] = input_vector[239] << 2;
assign MEM[1918] = input_vector[239] << 1;
assign MEM[1919] = input_vector[239] << 0;
assign MEM[1920] = -(input_vector[240] << 7);
assign MEM[1921] = input_vector[240] << 6;
assign MEM[1922] = input_vector[240] << 5;
assign MEM[1923] = input_vector[240] << 4;
assign MEM[1924] = input_vector[240] << 3;
assign MEM[1925] = input_vector[240] << 2;
assign MEM[1926] = input_vector[240] << 1;
assign MEM[1927] = input_vector[240] << 0;
assign MEM[1928] = -(input_vector[241] << 7);
assign MEM[1929] = input_vector[241] << 6;
assign MEM[1930] = input_vector[241] << 5;
assign MEM[1931] = input_vector[241] << 4;
assign MEM[1932] = input_vector[241] << 3;
assign MEM[1933] = input_vector[241] << 2;
assign MEM[1934] = input_vector[241] << 1;
assign MEM[1935] = input_vector[241] << 0;
assign MEM[1936] = -(input_vector[242] << 7);
assign MEM[1937] = input_vector[242] << 6;
assign MEM[1938] = input_vector[242] << 5;
assign MEM[1939] = input_vector[242] << 4;
assign MEM[1940] = input_vector[242] << 3;
assign MEM[1941] = input_vector[242] << 2;
assign MEM[1942] = input_vector[242] << 1;
assign MEM[1943] = input_vector[242] << 0;
assign MEM[1944] = -(input_vector[243] << 7);
assign MEM[1945] = input_vector[243] << 6;
assign MEM[1946] = input_vector[243] << 5;
assign MEM[1947] = input_vector[243] << 4;
assign MEM[1948] = input_vector[243] << 3;
assign MEM[1949] = input_vector[243] << 2;
assign MEM[1950] = input_vector[243] << 1;
assign MEM[1951] = input_vector[243] << 0;
assign MEM[1952] = -(input_vector[244] << 7);
assign MEM[1953] = input_vector[244] << 6;
assign MEM[1954] = input_vector[244] << 5;
assign MEM[1955] = input_vector[244] << 4;
assign MEM[1956] = input_vector[244] << 3;
assign MEM[1957] = input_vector[244] << 2;
assign MEM[1958] = input_vector[244] << 1;
assign MEM[1959] = input_vector[244] << 0;
assign MEM[1960] = -(input_vector[245] << 7);
assign MEM[1961] = input_vector[245] << 6;
assign MEM[1962] = input_vector[245] << 5;
assign MEM[1963] = input_vector[245] << 4;
assign MEM[1964] = input_vector[245] << 3;
assign MEM[1965] = input_vector[245] << 2;
assign MEM[1966] = input_vector[245] << 1;
assign MEM[1967] = input_vector[245] << 0;
assign MEM[1968] = -(input_vector[246] << 7);
assign MEM[1969] = input_vector[246] << 6;
assign MEM[1970] = input_vector[246] << 5;
assign MEM[1971] = input_vector[246] << 4;
assign MEM[1972] = input_vector[246] << 3;
assign MEM[1973] = input_vector[246] << 2;
assign MEM[1974] = input_vector[246] << 1;
assign MEM[1975] = input_vector[246] << 0;
assign MEM[1976] = -(input_vector[247] << 7);
assign MEM[1977] = input_vector[247] << 6;
assign MEM[1978] = input_vector[247] << 5;
assign MEM[1979] = input_vector[247] << 4;
assign MEM[1980] = input_vector[247] << 3;
assign MEM[1981] = input_vector[247] << 2;
assign MEM[1982] = input_vector[247] << 1;
assign MEM[1983] = input_vector[247] << 0;
assign MEM[1984] = -(input_vector[248] << 7);
assign MEM[1985] = input_vector[248] << 6;
assign MEM[1986] = input_vector[248] << 5;
assign MEM[1987] = input_vector[248] << 4;
assign MEM[1988] = input_vector[248] << 3;
assign MEM[1989] = input_vector[248] << 2;
assign MEM[1990] = input_vector[248] << 1;
assign MEM[1991] = input_vector[248] << 0;
assign MEM[1992] = -(input_vector[249] << 7);
assign MEM[1993] = input_vector[249] << 6;
assign MEM[1994] = input_vector[249] << 5;
assign MEM[1995] = input_vector[249] << 4;
assign MEM[1996] = input_vector[249] << 3;
assign MEM[1997] = input_vector[249] << 2;
assign MEM[1998] = input_vector[249] << 1;
assign MEM[1999] = input_vector[249] << 0;
assign MEM[2000] = -(input_vector[250] << 7);
assign MEM[2001] = input_vector[250] << 6;
assign MEM[2002] = input_vector[250] << 5;
assign MEM[2003] = input_vector[250] << 4;
assign MEM[2004] = input_vector[250] << 3;
assign MEM[2005] = input_vector[250] << 2;
assign MEM[2006] = input_vector[250] << 1;
assign MEM[2007] = input_vector[250] << 0;
assign MEM[2008] = -(input_vector[251] << 7);
assign MEM[2009] = input_vector[251] << 6;
assign MEM[2010] = input_vector[251] << 5;
assign MEM[2011] = input_vector[251] << 4;
assign MEM[2012] = input_vector[251] << 3;
assign MEM[2013] = input_vector[251] << 2;
assign MEM[2014] = input_vector[251] << 1;
assign MEM[2015] = input_vector[251] << 0;
assign MEM[2016] = -(input_vector[252] << 7);
assign MEM[2017] = input_vector[252] << 6;
assign MEM[2018] = input_vector[252] << 5;
assign MEM[2019] = input_vector[252] << 4;
assign MEM[2020] = input_vector[252] << 3;
assign MEM[2021] = input_vector[252] << 2;
assign MEM[2022] = input_vector[252] << 1;
assign MEM[2023] = input_vector[252] << 0;
assign MEM[2024] = -(input_vector[253] << 7);
assign MEM[2025] = input_vector[253] << 6;
assign MEM[2026] = input_vector[253] << 5;
assign MEM[2027] = input_vector[253] << 4;
assign MEM[2028] = input_vector[253] << 3;
assign MEM[2029] = input_vector[253] << 2;
assign MEM[2030] = input_vector[253] << 1;
assign MEM[2031] = input_vector[253] << 0;
assign MEM[2032] = -(input_vector[254] << 7);
assign MEM[2033] = input_vector[254] << 6;
assign MEM[2034] = input_vector[254] << 5;
assign MEM[2035] = input_vector[254] << 4;
assign MEM[2036] = input_vector[254] << 3;
assign MEM[2037] = input_vector[254] << 2;
assign MEM[2038] = input_vector[254] << 1;
assign MEM[2039] = input_vector[254] << 0;
assign MEM[2040] = -(input_vector[255] << 7);
assign MEM[2041] = input_vector[255] << 6;
assign MEM[2042] = input_vector[255] << 5;
assign MEM[2043] = input_vector[255] << 4;
assign MEM[2044] = input_vector[255] << 3;
assign MEM[2045] = input_vector[255] << 2;
assign MEM[2046] = input_vector[255] << 1;
assign MEM[2047] = input_vector[255] << 0;
assign MEM[2048] = -(input_vector[256] << 7);
assign MEM[2049] = input_vector[256] << 6;
assign MEM[2050] = input_vector[256] << 5;
assign MEM[2051] = input_vector[256] << 4;
assign MEM[2052] = input_vector[256] << 3;
assign MEM[2053] = input_vector[256] << 2;
assign MEM[2054] = input_vector[256] << 1;
assign MEM[2055] = input_vector[256] << 0;
assign MEM[2056] = -(input_vector[257] << 7);
assign MEM[2057] = input_vector[257] << 6;
assign MEM[2058] = input_vector[257] << 5;
assign MEM[2059] = input_vector[257] << 4;
assign MEM[2060] = input_vector[257] << 3;
assign MEM[2061] = input_vector[257] << 2;
assign MEM[2062] = input_vector[257] << 1;
assign MEM[2063] = input_vector[257] << 0;
assign MEM[2064] = -(input_vector[258] << 7);
assign MEM[2065] = input_vector[258] << 6;
assign MEM[2066] = input_vector[258] << 5;
assign MEM[2067] = input_vector[258] << 4;
assign MEM[2068] = input_vector[258] << 3;
assign MEM[2069] = input_vector[258] << 2;
assign MEM[2070] = input_vector[258] << 1;
assign MEM[2071] = input_vector[258] << 0;
assign MEM[2072] = -(input_vector[259] << 7);
assign MEM[2073] = input_vector[259] << 6;
assign MEM[2074] = input_vector[259] << 5;
assign MEM[2075] = input_vector[259] << 4;
assign MEM[2076] = input_vector[259] << 3;
assign MEM[2077] = input_vector[259] << 2;
assign MEM[2078] = input_vector[259] << 1;
assign MEM[2079] = input_vector[259] << 0;
assign MEM[2080] = -(input_vector[260] << 7);
assign MEM[2081] = input_vector[260] << 6;
assign MEM[2082] = input_vector[260] << 5;
assign MEM[2083] = input_vector[260] << 4;
assign MEM[2084] = input_vector[260] << 3;
assign MEM[2085] = input_vector[260] << 2;
assign MEM[2086] = input_vector[260] << 1;
assign MEM[2087] = input_vector[260] << 0;
assign MEM[2088] = -(input_vector[261] << 7);
assign MEM[2089] = input_vector[261] << 6;
assign MEM[2090] = input_vector[261] << 5;
assign MEM[2091] = input_vector[261] << 4;
assign MEM[2092] = input_vector[261] << 3;
assign MEM[2093] = input_vector[261] << 2;
assign MEM[2094] = input_vector[261] << 1;
assign MEM[2095] = input_vector[261] << 0;
assign MEM[2096] = -(input_vector[262] << 7);
assign MEM[2097] = input_vector[262] << 6;
assign MEM[2098] = input_vector[262] << 5;
assign MEM[2099] = input_vector[262] << 4;
assign MEM[2100] = input_vector[262] << 3;
assign MEM[2101] = input_vector[262] << 2;
assign MEM[2102] = input_vector[262] << 1;
assign MEM[2103] = input_vector[262] << 0;
assign MEM[2104] = -(input_vector[263] << 7);
assign MEM[2105] = input_vector[263] << 6;
assign MEM[2106] = input_vector[263] << 5;
assign MEM[2107] = input_vector[263] << 4;
assign MEM[2108] = input_vector[263] << 3;
assign MEM[2109] = input_vector[263] << 2;
assign MEM[2110] = input_vector[263] << 1;
assign MEM[2111] = input_vector[263] << 0;
assign MEM[2112] = -(input_vector[264] << 7);
assign MEM[2113] = input_vector[264] << 6;
assign MEM[2114] = input_vector[264] << 5;
assign MEM[2115] = input_vector[264] << 4;
assign MEM[2116] = input_vector[264] << 3;
assign MEM[2117] = input_vector[264] << 2;
assign MEM[2118] = input_vector[264] << 1;
assign MEM[2119] = input_vector[264] << 0;
assign MEM[2120] = -(input_vector[265] << 7);
assign MEM[2121] = input_vector[265] << 6;
assign MEM[2122] = input_vector[265] << 5;
assign MEM[2123] = input_vector[265] << 4;
assign MEM[2124] = input_vector[265] << 3;
assign MEM[2125] = input_vector[265] << 2;
assign MEM[2126] = input_vector[265] << 1;
assign MEM[2127] = input_vector[265] << 0;
assign MEM[2128] = -(input_vector[266] << 7);
assign MEM[2129] = input_vector[266] << 6;
assign MEM[2130] = input_vector[266] << 5;
assign MEM[2131] = input_vector[266] << 4;
assign MEM[2132] = input_vector[266] << 3;
assign MEM[2133] = input_vector[266] << 2;
assign MEM[2134] = input_vector[266] << 1;
assign MEM[2135] = input_vector[266] << 0;
assign MEM[2136] = -(input_vector[267] << 7);
assign MEM[2137] = input_vector[267] << 6;
assign MEM[2138] = input_vector[267] << 5;
assign MEM[2139] = input_vector[267] << 4;
assign MEM[2140] = input_vector[267] << 3;
assign MEM[2141] = input_vector[267] << 2;
assign MEM[2142] = input_vector[267] << 1;
assign MEM[2143] = input_vector[267] << 0;
assign MEM[2144] = -(input_vector[268] << 7);
assign MEM[2145] = input_vector[268] << 6;
assign MEM[2146] = input_vector[268] << 5;
assign MEM[2147] = input_vector[268] << 4;
assign MEM[2148] = input_vector[268] << 3;
assign MEM[2149] = input_vector[268] << 2;
assign MEM[2150] = input_vector[268] << 1;
assign MEM[2151] = input_vector[268] << 0;
assign MEM[2152] = -(input_vector[269] << 7);
assign MEM[2153] = input_vector[269] << 6;
assign MEM[2154] = input_vector[269] << 5;
assign MEM[2155] = input_vector[269] << 4;
assign MEM[2156] = input_vector[269] << 3;
assign MEM[2157] = input_vector[269] << 2;
assign MEM[2158] = input_vector[269] << 1;
assign MEM[2159] = input_vector[269] << 0;
assign MEM[2160] = -(input_vector[270] << 7);
assign MEM[2161] = input_vector[270] << 6;
assign MEM[2162] = input_vector[270] << 5;
assign MEM[2163] = input_vector[270] << 4;
assign MEM[2164] = input_vector[270] << 3;
assign MEM[2165] = input_vector[270] << 2;
assign MEM[2166] = input_vector[270] << 1;
assign MEM[2167] = input_vector[270] << 0;
assign MEM[2168] = -(input_vector[271] << 7);
assign MEM[2169] = input_vector[271] << 6;
assign MEM[2170] = input_vector[271] << 5;
assign MEM[2171] = input_vector[271] << 4;
assign MEM[2172] = input_vector[271] << 3;
assign MEM[2173] = input_vector[271] << 2;
assign MEM[2174] = input_vector[271] << 1;
assign MEM[2175] = input_vector[271] << 0;
assign MEM[2176] = -(input_vector[272] << 7);
assign MEM[2177] = input_vector[272] << 6;
assign MEM[2178] = input_vector[272] << 5;
assign MEM[2179] = input_vector[272] << 4;
assign MEM[2180] = input_vector[272] << 3;
assign MEM[2181] = input_vector[272] << 2;
assign MEM[2182] = input_vector[272] << 1;
assign MEM[2183] = input_vector[272] << 0;
assign MEM[2184] = -(input_vector[273] << 7);
assign MEM[2185] = input_vector[273] << 6;
assign MEM[2186] = input_vector[273] << 5;
assign MEM[2187] = input_vector[273] << 4;
assign MEM[2188] = input_vector[273] << 3;
assign MEM[2189] = input_vector[273] << 2;
assign MEM[2190] = input_vector[273] << 1;
assign MEM[2191] = input_vector[273] << 0;
assign MEM[2192] = -(input_vector[274] << 7);
assign MEM[2193] = input_vector[274] << 6;
assign MEM[2194] = input_vector[274] << 5;
assign MEM[2195] = input_vector[274] << 4;
assign MEM[2196] = input_vector[274] << 3;
assign MEM[2197] = input_vector[274] << 2;
assign MEM[2198] = input_vector[274] << 1;
assign MEM[2199] = input_vector[274] << 0;
assign MEM[2200] = -(input_vector[275] << 7);
assign MEM[2201] = input_vector[275] << 6;
assign MEM[2202] = input_vector[275] << 5;
assign MEM[2203] = input_vector[275] << 4;
assign MEM[2204] = input_vector[275] << 3;
assign MEM[2205] = input_vector[275] << 2;
assign MEM[2206] = input_vector[275] << 1;
assign MEM[2207] = input_vector[275] << 0;
assign MEM[2208] = -(input_vector[276] << 7);
assign MEM[2209] = input_vector[276] << 6;
assign MEM[2210] = input_vector[276] << 5;
assign MEM[2211] = input_vector[276] << 4;
assign MEM[2212] = input_vector[276] << 3;
assign MEM[2213] = input_vector[276] << 2;
assign MEM[2214] = input_vector[276] << 1;
assign MEM[2215] = input_vector[276] << 0;
assign MEM[2216] = -(input_vector[277] << 7);
assign MEM[2217] = input_vector[277] << 6;
assign MEM[2218] = input_vector[277] << 5;
assign MEM[2219] = input_vector[277] << 4;
assign MEM[2220] = input_vector[277] << 3;
assign MEM[2221] = input_vector[277] << 2;
assign MEM[2222] = input_vector[277] << 1;
assign MEM[2223] = input_vector[277] << 0;
assign MEM[2224] = -(input_vector[278] << 7);
assign MEM[2225] = input_vector[278] << 6;
assign MEM[2226] = input_vector[278] << 5;
assign MEM[2227] = input_vector[278] << 4;
assign MEM[2228] = input_vector[278] << 3;
assign MEM[2229] = input_vector[278] << 2;
assign MEM[2230] = input_vector[278] << 1;
assign MEM[2231] = input_vector[278] << 0;
assign MEM[2232] = -(input_vector[279] << 7);
assign MEM[2233] = input_vector[279] << 6;
assign MEM[2234] = input_vector[279] << 5;
assign MEM[2235] = input_vector[279] << 4;
assign MEM[2236] = input_vector[279] << 3;
assign MEM[2237] = input_vector[279] << 2;
assign MEM[2238] = input_vector[279] << 1;
assign MEM[2239] = input_vector[279] << 0;
assign MEM[2240] = -(input_vector[280] << 7);
assign MEM[2241] = input_vector[280] << 6;
assign MEM[2242] = input_vector[280] << 5;
assign MEM[2243] = input_vector[280] << 4;
assign MEM[2244] = input_vector[280] << 3;
assign MEM[2245] = input_vector[280] << 2;
assign MEM[2246] = input_vector[280] << 1;
assign MEM[2247] = input_vector[280] << 0;
assign MEM[2248] = -(input_vector[281] << 7);
assign MEM[2249] = input_vector[281] << 6;
assign MEM[2250] = input_vector[281] << 5;
assign MEM[2251] = input_vector[281] << 4;
assign MEM[2252] = input_vector[281] << 3;
assign MEM[2253] = input_vector[281] << 2;
assign MEM[2254] = input_vector[281] << 1;
assign MEM[2255] = input_vector[281] << 0;
assign MEM[2256] = -(input_vector[282] << 7);
assign MEM[2257] = input_vector[282] << 6;
assign MEM[2258] = input_vector[282] << 5;
assign MEM[2259] = input_vector[282] << 4;
assign MEM[2260] = input_vector[282] << 3;
assign MEM[2261] = input_vector[282] << 2;
assign MEM[2262] = input_vector[282] << 1;
assign MEM[2263] = input_vector[282] << 0;
assign MEM[2264] = -(input_vector[283] << 7);
assign MEM[2265] = input_vector[283] << 6;
assign MEM[2266] = input_vector[283] << 5;
assign MEM[2267] = input_vector[283] << 4;
assign MEM[2268] = input_vector[283] << 3;
assign MEM[2269] = input_vector[283] << 2;
assign MEM[2270] = input_vector[283] << 1;
assign MEM[2271] = input_vector[283] << 0;
assign MEM[2272] = -(input_vector[284] << 7);
assign MEM[2273] = input_vector[284] << 6;
assign MEM[2274] = input_vector[284] << 5;
assign MEM[2275] = input_vector[284] << 4;
assign MEM[2276] = input_vector[284] << 3;
assign MEM[2277] = input_vector[284] << 2;
assign MEM[2278] = input_vector[284] << 1;
assign MEM[2279] = input_vector[284] << 0;
assign MEM[2280] = -(input_vector[285] << 7);
assign MEM[2281] = input_vector[285] << 6;
assign MEM[2282] = input_vector[285] << 5;
assign MEM[2283] = input_vector[285] << 4;
assign MEM[2284] = input_vector[285] << 3;
assign MEM[2285] = input_vector[285] << 2;
assign MEM[2286] = input_vector[285] << 1;
assign MEM[2287] = input_vector[285] << 0;
assign MEM[2288] = -(input_vector[286] << 7);
assign MEM[2289] = input_vector[286] << 6;
assign MEM[2290] = input_vector[286] << 5;
assign MEM[2291] = input_vector[286] << 4;
assign MEM[2292] = input_vector[286] << 3;
assign MEM[2293] = input_vector[286] << 2;
assign MEM[2294] = input_vector[286] << 1;
assign MEM[2295] = input_vector[286] << 0;
assign MEM[2296] = -(input_vector[287] << 7);
assign MEM[2297] = input_vector[287] << 6;
assign MEM[2298] = input_vector[287] << 5;
assign MEM[2299] = input_vector[287] << 4;
assign MEM[2300] = input_vector[287] << 3;
assign MEM[2301] = input_vector[287] << 2;
assign MEM[2302] = input_vector[287] << 1;
assign MEM[2303] = input_vector[287] << 0;
assign MEM[2304] = -(input_vector[288] << 7);
assign MEM[2305] = input_vector[288] << 6;
assign MEM[2306] = input_vector[288] << 5;
assign MEM[2307] = input_vector[288] << 4;
assign MEM[2308] = input_vector[288] << 3;
assign MEM[2309] = input_vector[288] << 2;
assign MEM[2310] = input_vector[288] << 1;
assign MEM[2311] = input_vector[288] << 0;
assign MEM[2312] = -(input_vector[289] << 7);
assign MEM[2313] = input_vector[289] << 6;
assign MEM[2314] = input_vector[289] << 5;
assign MEM[2315] = input_vector[289] << 4;
assign MEM[2316] = input_vector[289] << 3;
assign MEM[2317] = input_vector[289] << 2;
assign MEM[2318] = input_vector[289] << 1;
assign MEM[2319] = input_vector[289] << 0;
assign MEM[2320] = -(input_vector[290] << 7);
assign MEM[2321] = input_vector[290] << 6;
assign MEM[2322] = input_vector[290] << 5;
assign MEM[2323] = input_vector[290] << 4;
assign MEM[2324] = input_vector[290] << 3;
assign MEM[2325] = input_vector[290] << 2;
assign MEM[2326] = input_vector[290] << 1;
assign MEM[2327] = input_vector[290] << 0;
assign MEM[2328] = -(input_vector[291] << 7);
assign MEM[2329] = input_vector[291] << 6;
assign MEM[2330] = input_vector[291] << 5;
assign MEM[2331] = input_vector[291] << 4;
assign MEM[2332] = input_vector[291] << 3;
assign MEM[2333] = input_vector[291] << 2;
assign MEM[2334] = input_vector[291] << 1;
assign MEM[2335] = input_vector[291] << 0;
assign MEM[2336] = -(input_vector[292] << 7);
assign MEM[2337] = input_vector[292] << 6;
assign MEM[2338] = input_vector[292] << 5;
assign MEM[2339] = input_vector[292] << 4;
assign MEM[2340] = input_vector[292] << 3;
assign MEM[2341] = input_vector[292] << 2;
assign MEM[2342] = input_vector[292] << 1;
assign MEM[2343] = input_vector[292] << 0;
assign MEM[2344] = -(input_vector[293] << 7);
assign MEM[2345] = input_vector[293] << 6;
assign MEM[2346] = input_vector[293] << 5;
assign MEM[2347] = input_vector[293] << 4;
assign MEM[2348] = input_vector[293] << 3;
assign MEM[2349] = input_vector[293] << 2;
assign MEM[2350] = input_vector[293] << 1;
assign MEM[2351] = input_vector[293] << 0;
assign MEM[2352] = -(input_vector[294] << 7);
assign MEM[2353] = input_vector[294] << 6;
assign MEM[2354] = input_vector[294] << 5;
assign MEM[2355] = input_vector[294] << 4;
assign MEM[2356] = input_vector[294] << 3;
assign MEM[2357] = input_vector[294] << 2;
assign MEM[2358] = input_vector[294] << 1;
assign MEM[2359] = input_vector[294] << 0;
assign MEM[2360] = -(input_vector[295] << 7);
assign MEM[2361] = input_vector[295] << 6;
assign MEM[2362] = input_vector[295] << 5;
assign MEM[2363] = input_vector[295] << 4;
assign MEM[2364] = input_vector[295] << 3;
assign MEM[2365] = input_vector[295] << 2;
assign MEM[2366] = input_vector[295] << 1;
assign MEM[2367] = input_vector[295] << 0;
assign MEM[2368] = -(input_vector[296] << 7);
assign MEM[2369] = input_vector[296] << 6;
assign MEM[2370] = input_vector[296] << 5;
assign MEM[2371] = input_vector[296] << 4;
assign MEM[2372] = input_vector[296] << 3;
assign MEM[2373] = input_vector[296] << 2;
assign MEM[2374] = input_vector[296] << 1;
assign MEM[2375] = input_vector[296] << 0;
assign MEM[2376] = -(input_vector[297] << 7);
assign MEM[2377] = input_vector[297] << 6;
assign MEM[2378] = input_vector[297] << 5;
assign MEM[2379] = input_vector[297] << 4;
assign MEM[2380] = input_vector[297] << 3;
assign MEM[2381] = input_vector[297] << 2;
assign MEM[2382] = input_vector[297] << 1;
assign MEM[2383] = input_vector[297] << 0;
assign MEM[2384] = -(input_vector[298] << 7);
assign MEM[2385] = input_vector[298] << 6;
assign MEM[2386] = input_vector[298] << 5;
assign MEM[2387] = input_vector[298] << 4;
assign MEM[2388] = input_vector[298] << 3;
assign MEM[2389] = input_vector[298] << 2;
assign MEM[2390] = input_vector[298] << 1;
assign MEM[2391] = input_vector[298] << 0;
assign MEM[2392] = -(input_vector[299] << 7);
assign MEM[2393] = input_vector[299] << 6;
assign MEM[2394] = input_vector[299] << 5;
assign MEM[2395] = input_vector[299] << 4;
assign MEM[2396] = input_vector[299] << 3;
assign MEM[2397] = input_vector[299] << 2;
assign MEM[2398] = input_vector[299] << 1;
assign MEM[2399] = input_vector[299] << 0;
assign MEM[2400] = -(input_vector[300] << 7);
assign MEM[2401] = input_vector[300] << 6;
assign MEM[2402] = input_vector[300] << 5;
assign MEM[2403] = input_vector[300] << 4;
assign MEM[2404] = input_vector[300] << 3;
assign MEM[2405] = input_vector[300] << 2;
assign MEM[2406] = input_vector[300] << 1;
assign MEM[2407] = input_vector[300] << 0;
assign MEM[2408] = -(input_vector[301] << 7);
assign MEM[2409] = input_vector[301] << 6;
assign MEM[2410] = input_vector[301] << 5;
assign MEM[2411] = input_vector[301] << 4;
assign MEM[2412] = input_vector[301] << 3;
assign MEM[2413] = input_vector[301] << 2;
assign MEM[2414] = input_vector[301] << 1;
assign MEM[2415] = input_vector[301] << 0;
assign MEM[2416] = -(input_vector[302] << 7);
assign MEM[2417] = input_vector[302] << 6;
assign MEM[2418] = input_vector[302] << 5;
assign MEM[2419] = input_vector[302] << 4;
assign MEM[2420] = input_vector[302] << 3;
assign MEM[2421] = input_vector[302] << 2;
assign MEM[2422] = input_vector[302] << 1;
assign MEM[2423] = input_vector[302] << 0;
assign MEM[2424] = -(input_vector[303] << 7);
assign MEM[2425] = input_vector[303] << 6;
assign MEM[2426] = input_vector[303] << 5;
assign MEM[2427] = input_vector[303] << 4;
assign MEM[2428] = input_vector[303] << 3;
assign MEM[2429] = input_vector[303] << 2;
assign MEM[2430] = input_vector[303] << 1;
assign MEM[2431] = input_vector[303] << 0;
assign MEM[2432] = -(input_vector[304] << 7);
assign MEM[2433] = input_vector[304] << 6;
assign MEM[2434] = input_vector[304] << 5;
assign MEM[2435] = input_vector[304] << 4;
assign MEM[2436] = input_vector[304] << 3;
assign MEM[2437] = input_vector[304] << 2;
assign MEM[2438] = input_vector[304] << 1;
assign MEM[2439] = input_vector[304] << 0;
assign MEM[2440] = -(input_vector[305] << 7);
assign MEM[2441] = input_vector[305] << 6;
assign MEM[2442] = input_vector[305] << 5;
assign MEM[2443] = input_vector[305] << 4;
assign MEM[2444] = input_vector[305] << 3;
assign MEM[2445] = input_vector[305] << 2;
assign MEM[2446] = input_vector[305] << 1;
assign MEM[2447] = input_vector[305] << 0;
assign MEM[2448] = -(input_vector[306] << 7);
assign MEM[2449] = input_vector[306] << 6;
assign MEM[2450] = input_vector[306] << 5;
assign MEM[2451] = input_vector[306] << 4;
assign MEM[2452] = input_vector[306] << 3;
assign MEM[2453] = input_vector[306] << 2;
assign MEM[2454] = input_vector[306] << 1;
assign MEM[2455] = input_vector[306] << 0;
assign MEM[2456] = -(input_vector[307] << 7);
assign MEM[2457] = input_vector[307] << 6;
assign MEM[2458] = input_vector[307] << 5;
assign MEM[2459] = input_vector[307] << 4;
assign MEM[2460] = input_vector[307] << 3;
assign MEM[2461] = input_vector[307] << 2;
assign MEM[2462] = input_vector[307] << 1;
assign MEM[2463] = input_vector[307] << 0;
assign MEM[2464] = -(input_vector[308] << 7);
assign MEM[2465] = input_vector[308] << 6;
assign MEM[2466] = input_vector[308] << 5;
assign MEM[2467] = input_vector[308] << 4;
assign MEM[2468] = input_vector[308] << 3;
assign MEM[2469] = input_vector[308] << 2;
assign MEM[2470] = input_vector[308] << 1;
assign MEM[2471] = input_vector[308] << 0;
assign MEM[2472] = -(input_vector[309] << 7);
assign MEM[2473] = input_vector[309] << 6;
assign MEM[2474] = input_vector[309] << 5;
assign MEM[2475] = input_vector[309] << 4;
assign MEM[2476] = input_vector[309] << 3;
assign MEM[2477] = input_vector[309] << 2;
assign MEM[2478] = input_vector[309] << 1;
assign MEM[2479] = input_vector[309] << 0;
assign MEM[2480] = -(input_vector[310] << 7);
assign MEM[2481] = input_vector[310] << 6;
assign MEM[2482] = input_vector[310] << 5;
assign MEM[2483] = input_vector[310] << 4;
assign MEM[2484] = input_vector[310] << 3;
assign MEM[2485] = input_vector[310] << 2;
assign MEM[2486] = input_vector[310] << 1;
assign MEM[2487] = input_vector[310] << 0;
assign MEM[2488] = -(input_vector[311] << 7);
assign MEM[2489] = input_vector[311] << 6;
assign MEM[2490] = input_vector[311] << 5;
assign MEM[2491] = input_vector[311] << 4;
assign MEM[2492] = input_vector[311] << 3;
assign MEM[2493] = input_vector[311] << 2;
assign MEM[2494] = input_vector[311] << 1;
assign MEM[2495] = input_vector[311] << 0;
assign MEM[2496] = -(input_vector[312] << 7);
assign MEM[2497] = input_vector[312] << 6;
assign MEM[2498] = input_vector[312] << 5;
assign MEM[2499] = input_vector[312] << 4;
assign MEM[2500] = input_vector[312] << 3;
assign MEM[2501] = input_vector[312] << 2;
assign MEM[2502] = input_vector[312] << 1;
assign MEM[2503] = input_vector[312] << 0;
assign MEM[2504] = -(input_vector[313] << 7);
assign MEM[2505] = input_vector[313] << 6;
assign MEM[2506] = input_vector[313] << 5;
assign MEM[2507] = input_vector[313] << 4;
assign MEM[2508] = input_vector[313] << 3;
assign MEM[2509] = input_vector[313] << 2;
assign MEM[2510] = input_vector[313] << 1;
assign MEM[2511] = input_vector[313] << 0;
assign MEM[2512] = -(input_vector[314] << 7);
assign MEM[2513] = input_vector[314] << 6;
assign MEM[2514] = input_vector[314] << 5;
assign MEM[2515] = input_vector[314] << 4;
assign MEM[2516] = input_vector[314] << 3;
assign MEM[2517] = input_vector[314] << 2;
assign MEM[2518] = input_vector[314] << 1;
assign MEM[2519] = input_vector[314] << 0;
assign MEM[2520] = -(input_vector[315] << 7);
assign MEM[2521] = input_vector[315] << 6;
assign MEM[2522] = input_vector[315] << 5;
assign MEM[2523] = input_vector[315] << 4;
assign MEM[2524] = input_vector[315] << 3;
assign MEM[2525] = input_vector[315] << 2;
assign MEM[2526] = input_vector[315] << 1;
assign MEM[2527] = input_vector[315] << 0;
assign MEM[2528] = -(input_vector[316] << 7);
assign MEM[2529] = input_vector[316] << 6;
assign MEM[2530] = input_vector[316] << 5;
assign MEM[2531] = input_vector[316] << 4;
assign MEM[2532] = input_vector[316] << 3;
assign MEM[2533] = input_vector[316] << 2;
assign MEM[2534] = input_vector[316] << 1;
assign MEM[2535] = input_vector[316] << 0;
assign MEM[2536] = -(input_vector[317] << 7);
assign MEM[2537] = input_vector[317] << 6;
assign MEM[2538] = input_vector[317] << 5;
assign MEM[2539] = input_vector[317] << 4;
assign MEM[2540] = input_vector[317] << 3;
assign MEM[2541] = input_vector[317] << 2;
assign MEM[2542] = input_vector[317] << 1;
assign MEM[2543] = input_vector[317] << 0;
assign MEM[2544] = -(input_vector[318] << 7);
assign MEM[2545] = input_vector[318] << 6;
assign MEM[2546] = input_vector[318] << 5;
assign MEM[2547] = input_vector[318] << 4;
assign MEM[2548] = input_vector[318] << 3;
assign MEM[2549] = input_vector[318] << 2;
assign MEM[2550] = input_vector[318] << 1;
assign MEM[2551] = input_vector[318] << 0;
assign MEM[2552] = -(input_vector[319] << 7);
assign MEM[2553] = input_vector[319] << 6;
assign MEM[2554] = input_vector[319] << 5;
assign MEM[2555] = input_vector[319] << 4;
assign MEM[2556] = input_vector[319] << 3;
assign MEM[2557] = input_vector[319] << 2;
assign MEM[2558] = input_vector[319] << 1;
assign MEM[2559] = input_vector[319] << 0;
assign MEM[2560] = -(input_vector[320] << 7);
assign MEM[2561] = input_vector[320] << 6;
assign MEM[2562] = input_vector[320] << 5;
assign MEM[2563] = input_vector[320] << 4;
assign MEM[2564] = input_vector[320] << 3;
assign MEM[2565] = input_vector[320] << 2;
assign MEM[2566] = input_vector[320] << 1;
assign MEM[2567] = input_vector[320] << 0;
assign MEM[2568] = -(input_vector[321] << 7);
assign MEM[2569] = input_vector[321] << 6;
assign MEM[2570] = input_vector[321] << 5;
assign MEM[2571] = input_vector[321] << 4;
assign MEM[2572] = input_vector[321] << 3;
assign MEM[2573] = input_vector[321] << 2;
assign MEM[2574] = input_vector[321] << 1;
assign MEM[2575] = input_vector[321] << 0;
assign MEM[2576] = -(input_vector[322] << 7);
assign MEM[2577] = input_vector[322] << 6;
assign MEM[2578] = input_vector[322] << 5;
assign MEM[2579] = input_vector[322] << 4;
assign MEM[2580] = input_vector[322] << 3;
assign MEM[2581] = input_vector[322] << 2;
assign MEM[2582] = input_vector[322] << 1;
assign MEM[2583] = input_vector[322] << 0;
assign MEM[2584] = -(input_vector[323] << 7);
assign MEM[2585] = input_vector[323] << 6;
assign MEM[2586] = input_vector[323] << 5;
assign MEM[2587] = input_vector[323] << 4;
assign MEM[2588] = input_vector[323] << 3;
assign MEM[2589] = input_vector[323] << 2;
assign MEM[2590] = input_vector[323] << 1;
assign MEM[2591] = input_vector[323] << 0;
assign MEM[2592] = -(input_vector[324] << 7);
assign MEM[2593] = input_vector[324] << 6;
assign MEM[2594] = input_vector[324] << 5;
assign MEM[2595] = input_vector[324] << 4;
assign MEM[2596] = input_vector[324] << 3;
assign MEM[2597] = input_vector[324] << 2;
assign MEM[2598] = input_vector[324] << 1;
assign MEM[2599] = input_vector[324] << 0;
assign MEM[2600] = -(input_vector[325] << 7);
assign MEM[2601] = input_vector[325] << 6;
assign MEM[2602] = input_vector[325] << 5;
assign MEM[2603] = input_vector[325] << 4;
assign MEM[2604] = input_vector[325] << 3;
assign MEM[2605] = input_vector[325] << 2;
assign MEM[2606] = input_vector[325] << 1;
assign MEM[2607] = input_vector[325] << 0;
assign MEM[2608] = -(input_vector[326] << 7);
assign MEM[2609] = input_vector[326] << 6;
assign MEM[2610] = input_vector[326] << 5;
assign MEM[2611] = input_vector[326] << 4;
assign MEM[2612] = input_vector[326] << 3;
assign MEM[2613] = input_vector[326] << 2;
assign MEM[2614] = input_vector[326] << 1;
assign MEM[2615] = input_vector[326] << 0;
assign MEM[2616] = -(input_vector[327] << 7);
assign MEM[2617] = input_vector[327] << 6;
assign MEM[2618] = input_vector[327] << 5;
assign MEM[2619] = input_vector[327] << 4;
assign MEM[2620] = input_vector[327] << 3;
assign MEM[2621] = input_vector[327] << 2;
assign MEM[2622] = input_vector[327] << 1;
assign MEM[2623] = input_vector[327] << 0;
assign MEM[2624] = -(input_vector[328] << 7);
assign MEM[2625] = input_vector[328] << 6;
assign MEM[2626] = input_vector[328] << 5;
assign MEM[2627] = input_vector[328] << 4;
assign MEM[2628] = input_vector[328] << 3;
assign MEM[2629] = input_vector[328] << 2;
assign MEM[2630] = input_vector[328] << 1;
assign MEM[2631] = input_vector[328] << 0;
assign MEM[2632] = -(input_vector[329] << 7);
assign MEM[2633] = input_vector[329] << 6;
assign MEM[2634] = input_vector[329] << 5;
assign MEM[2635] = input_vector[329] << 4;
assign MEM[2636] = input_vector[329] << 3;
assign MEM[2637] = input_vector[329] << 2;
assign MEM[2638] = input_vector[329] << 1;
assign MEM[2639] = input_vector[329] << 0;
assign MEM[2640] = -(input_vector[330] << 7);
assign MEM[2641] = input_vector[330] << 6;
assign MEM[2642] = input_vector[330] << 5;
assign MEM[2643] = input_vector[330] << 4;
assign MEM[2644] = input_vector[330] << 3;
assign MEM[2645] = input_vector[330] << 2;
assign MEM[2646] = input_vector[330] << 1;
assign MEM[2647] = input_vector[330] << 0;
assign MEM[2648] = -(input_vector[331] << 7);
assign MEM[2649] = input_vector[331] << 6;
assign MEM[2650] = input_vector[331] << 5;
assign MEM[2651] = input_vector[331] << 4;
assign MEM[2652] = input_vector[331] << 3;
assign MEM[2653] = input_vector[331] << 2;
assign MEM[2654] = input_vector[331] << 1;
assign MEM[2655] = input_vector[331] << 0;
assign MEM[2656] = -(input_vector[332] << 7);
assign MEM[2657] = input_vector[332] << 6;
assign MEM[2658] = input_vector[332] << 5;
assign MEM[2659] = input_vector[332] << 4;
assign MEM[2660] = input_vector[332] << 3;
assign MEM[2661] = input_vector[332] << 2;
assign MEM[2662] = input_vector[332] << 1;
assign MEM[2663] = input_vector[332] << 0;
assign MEM[2664] = -(input_vector[333] << 7);
assign MEM[2665] = input_vector[333] << 6;
assign MEM[2666] = input_vector[333] << 5;
assign MEM[2667] = input_vector[333] << 4;
assign MEM[2668] = input_vector[333] << 3;
assign MEM[2669] = input_vector[333] << 2;
assign MEM[2670] = input_vector[333] << 1;
assign MEM[2671] = input_vector[333] << 0;
assign MEM[2672] = -(input_vector[334] << 7);
assign MEM[2673] = input_vector[334] << 6;
assign MEM[2674] = input_vector[334] << 5;
assign MEM[2675] = input_vector[334] << 4;
assign MEM[2676] = input_vector[334] << 3;
assign MEM[2677] = input_vector[334] << 2;
assign MEM[2678] = input_vector[334] << 1;
assign MEM[2679] = input_vector[334] << 0;
assign MEM[2680] = -(input_vector[335] << 7);
assign MEM[2681] = input_vector[335] << 6;
assign MEM[2682] = input_vector[335] << 5;
assign MEM[2683] = input_vector[335] << 4;
assign MEM[2684] = input_vector[335] << 3;
assign MEM[2685] = input_vector[335] << 2;
assign MEM[2686] = input_vector[335] << 1;
assign MEM[2687] = input_vector[335] << 0;
assign MEM[2688] = -(input_vector[336] << 7);
assign MEM[2689] = input_vector[336] << 6;
assign MEM[2690] = input_vector[336] << 5;
assign MEM[2691] = input_vector[336] << 4;
assign MEM[2692] = input_vector[336] << 3;
assign MEM[2693] = input_vector[336] << 2;
assign MEM[2694] = input_vector[336] << 1;
assign MEM[2695] = input_vector[336] << 0;
assign MEM[2696] = -(input_vector[337] << 7);
assign MEM[2697] = input_vector[337] << 6;
assign MEM[2698] = input_vector[337] << 5;
assign MEM[2699] = input_vector[337] << 4;
assign MEM[2700] = input_vector[337] << 3;
assign MEM[2701] = input_vector[337] << 2;
assign MEM[2702] = input_vector[337] << 1;
assign MEM[2703] = input_vector[337] << 0;
assign MEM[2704] = -(input_vector[338] << 7);
assign MEM[2705] = input_vector[338] << 6;
assign MEM[2706] = input_vector[338] << 5;
assign MEM[2707] = input_vector[338] << 4;
assign MEM[2708] = input_vector[338] << 3;
assign MEM[2709] = input_vector[338] << 2;
assign MEM[2710] = input_vector[338] << 1;
assign MEM[2711] = input_vector[338] << 0;
assign MEM[2712] = -(input_vector[339] << 7);
assign MEM[2713] = input_vector[339] << 6;
assign MEM[2714] = input_vector[339] << 5;
assign MEM[2715] = input_vector[339] << 4;
assign MEM[2716] = input_vector[339] << 3;
assign MEM[2717] = input_vector[339] << 2;
assign MEM[2718] = input_vector[339] << 1;
assign MEM[2719] = input_vector[339] << 0;
assign MEM[2720] = -(input_vector[340] << 7);
assign MEM[2721] = input_vector[340] << 6;
assign MEM[2722] = input_vector[340] << 5;
assign MEM[2723] = input_vector[340] << 4;
assign MEM[2724] = input_vector[340] << 3;
assign MEM[2725] = input_vector[340] << 2;
assign MEM[2726] = input_vector[340] << 1;
assign MEM[2727] = input_vector[340] << 0;
assign MEM[2728] = -(input_vector[341] << 7);
assign MEM[2729] = input_vector[341] << 6;
assign MEM[2730] = input_vector[341] << 5;
assign MEM[2731] = input_vector[341] << 4;
assign MEM[2732] = input_vector[341] << 3;
assign MEM[2733] = input_vector[341] << 2;
assign MEM[2734] = input_vector[341] << 1;
assign MEM[2735] = input_vector[341] << 0;
assign MEM[2736] = -(input_vector[342] << 7);
assign MEM[2737] = input_vector[342] << 6;
assign MEM[2738] = input_vector[342] << 5;
assign MEM[2739] = input_vector[342] << 4;
assign MEM[2740] = input_vector[342] << 3;
assign MEM[2741] = input_vector[342] << 2;
assign MEM[2742] = input_vector[342] << 1;
assign MEM[2743] = input_vector[342] << 0;
assign MEM[2744] = -(input_vector[343] << 7);
assign MEM[2745] = input_vector[343] << 6;
assign MEM[2746] = input_vector[343] << 5;
assign MEM[2747] = input_vector[343] << 4;
assign MEM[2748] = input_vector[343] << 3;
assign MEM[2749] = input_vector[343] << 2;
assign MEM[2750] = input_vector[343] << 1;
assign MEM[2751] = input_vector[343] << 0;
assign MEM[2752] = -(input_vector[344] << 7);
assign MEM[2753] = input_vector[344] << 6;
assign MEM[2754] = input_vector[344] << 5;
assign MEM[2755] = input_vector[344] << 4;
assign MEM[2756] = input_vector[344] << 3;
assign MEM[2757] = input_vector[344] << 2;
assign MEM[2758] = input_vector[344] << 1;
assign MEM[2759] = input_vector[344] << 0;
assign MEM[2760] = -(input_vector[345] << 7);
assign MEM[2761] = input_vector[345] << 6;
assign MEM[2762] = input_vector[345] << 5;
assign MEM[2763] = input_vector[345] << 4;
assign MEM[2764] = input_vector[345] << 3;
assign MEM[2765] = input_vector[345] << 2;
assign MEM[2766] = input_vector[345] << 1;
assign MEM[2767] = input_vector[345] << 0;
assign MEM[2768] = -(input_vector[346] << 7);
assign MEM[2769] = input_vector[346] << 6;
assign MEM[2770] = input_vector[346] << 5;
assign MEM[2771] = input_vector[346] << 4;
assign MEM[2772] = input_vector[346] << 3;
assign MEM[2773] = input_vector[346] << 2;
assign MEM[2774] = input_vector[346] << 1;
assign MEM[2775] = input_vector[346] << 0;
assign MEM[2776] = -(input_vector[347] << 7);
assign MEM[2777] = input_vector[347] << 6;
assign MEM[2778] = input_vector[347] << 5;
assign MEM[2779] = input_vector[347] << 4;
assign MEM[2780] = input_vector[347] << 3;
assign MEM[2781] = input_vector[347] << 2;
assign MEM[2782] = input_vector[347] << 1;
assign MEM[2783] = input_vector[347] << 0;
assign MEM[2784] = -(input_vector[348] << 7);
assign MEM[2785] = input_vector[348] << 6;
assign MEM[2786] = input_vector[348] << 5;
assign MEM[2787] = input_vector[348] << 4;
assign MEM[2788] = input_vector[348] << 3;
assign MEM[2789] = input_vector[348] << 2;
assign MEM[2790] = input_vector[348] << 1;
assign MEM[2791] = input_vector[348] << 0;
assign MEM[2792] = -(input_vector[349] << 7);
assign MEM[2793] = input_vector[349] << 6;
assign MEM[2794] = input_vector[349] << 5;
assign MEM[2795] = input_vector[349] << 4;
assign MEM[2796] = input_vector[349] << 3;
assign MEM[2797] = input_vector[349] << 2;
assign MEM[2798] = input_vector[349] << 1;
assign MEM[2799] = input_vector[349] << 0;
assign MEM[2800] = -(input_vector[350] << 7);
assign MEM[2801] = input_vector[350] << 6;
assign MEM[2802] = input_vector[350] << 5;
assign MEM[2803] = input_vector[350] << 4;
assign MEM[2804] = input_vector[350] << 3;
assign MEM[2805] = input_vector[350] << 2;
assign MEM[2806] = input_vector[350] << 1;
assign MEM[2807] = input_vector[350] << 0;
assign MEM[2808] = -(input_vector[351] << 7);
assign MEM[2809] = input_vector[351] << 6;
assign MEM[2810] = input_vector[351] << 5;
assign MEM[2811] = input_vector[351] << 4;
assign MEM[2812] = input_vector[351] << 3;
assign MEM[2813] = input_vector[351] << 2;
assign MEM[2814] = input_vector[351] << 1;
assign MEM[2815] = input_vector[351] << 0;
assign MEM[2816] = -(input_vector[352] << 7);
assign MEM[2817] = input_vector[352] << 6;
assign MEM[2818] = input_vector[352] << 5;
assign MEM[2819] = input_vector[352] << 4;
assign MEM[2820] = input_vector[352] << 3;
assign MEM[2821] = input_vector[352] << 2;
assign MEM[2822] = input_vector[352] << 1;
assign MEM[2823] = input_vector[352] << 0;
assign MEM[2824] = -(input_vector[353] << 7);
assign MEM[2825] = input_vector[353] << 6;
assign MEM[2826] = input_vector[353] << 5;
assign MEM[2827] = input_vector[353] << 4;
assign MEM[2828] = input_vector[353] << 3;
assign MEM[2829] = input_vector[353] << 2;
assign MEM[2830] = input_vector[353] << 1;
assign MEM[2831] = input_vector[353] << 0;
assign MEM[2832] = -(input_vector[354] << 7);
assign MEM[2833] = input_vector[354] << 6;
assign MEM[2834] = input_vector[354] << 5;
assign MEM[2835] = input_vector[354] << 4;
assign MEM[2836] = input_vector[354] << 3;
assign MEM[2837] = input_vector[354] << 2;
assign MEM[2838] = input_vector[354] << 1;
assign MEM[2839] = input_vector[354] << 0;
assign MEM[2840] = -(input_vector[355] << 7);
assign MEM[2841] = input_vector[355] << 6;
assign MEM[2842] = input_vector[355] << 5;
assign MEM[2843] = input_vector[355] << 4;
assign MEM[2844] = input_vector[355] << 3;
assign MEM[2845] = input_vector[355] << 2;
assign MEM[2846] = input_vector[355] << 1;
assign MEM[2847] = input_vector[355] << 0;
assign MEM[2848] = -(input_vector[356] << 7);
assign MEM[2849] = input_vector[356] << 6;
assign MEM[2850] = input_vector[356] << 5;
assign MEM[2851] = input_vector[356] << 4;
assign MEM[2852] = input_vector[356] << 3;
assign MEM[2853] = input_vector[356] << 2;
assign MEM[2854] = input_vector[356] << 1;
assign MEM[2855] = input_vector[356] << 0;
assign MEM[2856] = -(input_vector[357] << 7);
assign MEM[2857] = input_vector[357] << 6;
assign MEM[2858] = input_vector[357] << 5;
assign MEM[2859] = input_vector[357] << 4;
assign MEM[2860] = input_vector[357] << 3;
assign MEM[2861] = input_vector[357] << 2;
assign MEM[2862] = input_vector[357] << 1;
assign MEM[2863] = input_vector[357] << 0;
assign MEM[2864] = -(input_vector[358] << 7);
assign MEM[2865] = input_vector[358] << 6;
assign MEM[2866] = input_vector[358] << 5;
assign MEM[2867] = input_vector[358] << 4;
assign MEM[2868] = input_vector[358] << 3;
assign MEM[2869] = input_vector[358] << 2;
assign MEM[2870] = input_vector[358] << 1;
assign MEM[2871] = input_vector[358] << 0;
assign MEM[2872] = -(input_vector[359] << 7);
assign MEM[2873] = input_vector[359] << 6;
assign MEM[2874] = input_vector[359] << 5;
assign MEM[2875] = input_vector[359] << 4;
assign MEM[2876] = input_vector[359] << 3;
assign MEM[2877] = input_vector[359] << 2;
assign MEM[2878] = input_vector[359] << 1;
assign MEM[2879] = input_vector[359] << 0;
assign MEM[2880] = -(input_vector[360] << 7);
assign MEM[2881] = input_vector[360] << 6;
assign MEM[2882] = input_vector[360] << 5;
assign MEM[2883] = input_vector[360] << 4;
assign MEM[2884] = input_vector[360] << 3;
assign MEM[2885] = input_vector[360] << 2;
assign MEM[2886] = input_vector[360] << 1;
assign MEM[2887] = input_vector[360] << 0;
assign MEM[2888] = -(input_vector[361] << 7);
assign MEM[2889] = input_vector[361] << 6;
assign MEM[2890] = input_vector[361] << 5;
assign MEM[2891] = input_vector[361] << 4;
assign MEM[2892] = input_vector[361] << 3;
assign MEM[2893] = input_vector[361] << 2;
assign MEM[2894] = input_vector[361] << 1;
assign MEM[2895] = input_vector[361] << 0;
assign MEM[2896] = -(input_vector[362] << 7);
assign MEM[2897] = input_vector[362] << 6;
assign MEM[2898] = input_vector[362] << 5;
assign MEM[2899] = input_vector[362] << 4;
assign MEM[2900] = input_vector[362] << 3;
assign MEM[2901] = input_vector[362] << 2;
assign MEM[2902] = input_vector[362] << 1;
assign MEM[2903] = input_vector[362] << 0;
assign MEM[2904] = -(input_vector[363] << 7);
assign MEM[2905] = input_vector[363] << 6;
assign MEM[2906] = input_vector[363] << 5;
assign MEM[2907] = input_vector[363] << 4;
assign MEM[2908] = input_vector[363] << 3;
assign MEM[2909] = input_vector[363] << 2;
assign MEM[2910] = input_vector[363] << 1;
assign MEM[2911] = input_vector[363] << 0;
assign MEM[2912] = -(input_vector[364] << 7);
assign MEM[2913] = input_vector[364] << 6;
assign MEM[2914] = input_vector[364] << 5;
assign MEM[2915] = input_vector[364] << 4;
assign MEM[2916] = input_vector[364] << 3;
assign MEM[2917] = input_vector[364] << 2;
assign MEM[2918] = input_vector[364] << 1;
assign MEM[2919] = input_vector[364] << 0;
assign MEM[2920] = -(input_vector[365] << 7);
assign MEM[2921] = input_vector[365] << 6;
assign MEM[2922] = input_vector[365] << 5;
assign MEM[2923] = input_vector[365] << 4;
assign MEM[2924] = input_vector[365] << 3;
assign MEM[2925] = input_vector[365] << 2;
assign MEM[2926] = input_vector[365] << 1;
assign MEM[2927] = input_vector[365] << 0;
assign MEM[2928] = -(input_vector[366] << 7);
assign MEM[2929] = input_vector[366] << 6;
assign MEM[2930] = input_vector[366] << 5;
assign MEM[2931] = input_vector[366] << 4;
assign MEM[2932] = input_vector[366] << 3;
assign MEM[2933] = input_vector[366] << 2;
assign MEM[2934] = input_vector[366] << 1;
assign MEM[2935] = input_vector[366] << 0;
assign MEM[2936] = -(input_vector[367] << 7);
assign MEM[2937] = input_vector[367] << 6;
assign MEM[2938] = input_vector[367] << 5;
assign MEM[2939] = input_vector[367] << 4;
assign MEM[2940] = input_vector[367] << 3;
assign MEM[2941] = input_vector[367] << 2;
assign MEM[2942] = input_vector[367] << 1;
assign MEM[2943] = input_vector[367] << 0;
assign MEM[2944] = -(input_vector[368] << 7);
assign MEM[2945] = input_vector[368] << 6;
assign MEM[2946] = input_vector[368] << 5;
assign MEM[2947] = input_vector[368] << 4;
assign MEM[2948] = input_vector[368] << 3;
assign MEM[2949] = input_vector[368] << 2;
assign MEM[2950] = input_vector[368] << 1;
assign MEM[2951] = input_vector[368] << 0;
assign MEM[2952] = -(input_vector[369] << 7);
assign MEM[2953] = input_vector[369] << 6;
assign MEM[2954] = input_vector[369] << 5;
assign MEM[2955] = input_vector[369] << 4;
assign MEM[2956] = input_vector[369] << 3;
assign MEM[2957] = input_vector[369] << 2;
assign MEM[2958] = input_vector[369] << 1;
assign MEM[2959] = input_vector[369] << 0;
assign MEM[2960] = -(input_vector[370] << 7);
assign MEM[2961] = input_vector[370] << 6;
assign MEM[2962] = input_vector[370] << 5;
assign MEM[2963] = input_vector[370] << 4;
assign MEM[2964] = input_vector[370] << 3;
assign MEM[2965] = input_vector[370] << 2;
assign MEM[2966] = input_vector[370] << 1;
assign MEM[2967] = input_vector[370] << 0;
assign MEM[2968] = -(input_vector[371] << 7);
assign MEM[2969] = input_vector[371] << 6;
assign MEM[2970] = input_vector[371] << 5;
assign MEM[2971] = input_vector[371] << 4;
assign MEM[2972] = input_vector[371] << 3;
assign MEM[2973] = input_vector[371] << 2;
assign MEM[2974] = input_vector[371] << 1;
assign MEM[2975] = input_vector[371] << 0;
assign MEM[2976] = -(input_vector[372] << 7);
assign MEM[2977] = input_vector[372] << 6;
assign MEM[2978] = input_vector[372] << 5;
assign MEM[2979] = input_vector[372] << 4;
assign MEM[2980] = input_vector[372] << 3;
assign MEM[2981] = input_vector[372] << 2;
assign MEM[2982] = input_vector[372] << 1;
assign MEM[2983] = input_vector[372] << 0;
assign MEM[2984] = -(input_vector[373] << 7);
assign MEM[2985] = input_vector[373] << 6;
assign MEM[2986] = input_vector[373] << 5;
assign MEM[2987] = input_vector[373] << 4;
assign MEM[2988] = input_vector[373] << 3;
assign MEM[2989] = input_vector[373] << 2;
assign MEM[2990] = input_vector[373] << 1;
assign MEM[2991] = input_vector[373] << 0;
assign MEM[2992] = -(input_vector[374] << 7);
assign MEM[2993] = input_vector[374] << 6;
assign MEM[2994] = input_vector[374] << 5;
assign MEM[2995] = input_vector[374] << 4;
assign MEM[2996] = input_vector[374] << 3;
assign MEM[2997] = input_vector[374] << 2;
assign MEM[2998] = input_vector[374] << 1;
assign MEM[2999] = input_vector[374] << 0;
assign MEM[3000] = -(input_vector[375] << 7);
assign MEM[3001] = input_vector[375] << 6;
assign MEM[3002] = input_vector[375] << 5;
assign MEM[3003] = input_vector[375] << 4;
assign MEM[3004] = input_vector[375] << 3;
assign MEM[3005] = input_vector[375] << 2;
assign MEM[3006] = input_vector[375] << 1;
assign MEM[3007] = input_vector[375] << 0;
assign MEM[3008] = -(input_vector[376] << 7);
assign MEM[3009] = input_vector[376] << 6;
assign MEM[3010] = input_vector[376] << 5;
assign MEM[3011] = input_vector[376] << 4;
assign MEM[3012] = input_vector[376] << 3;
assign MEM[3013] = input_vector[376] << 2;
assign MEM[3014] = input_vector[376] << 1;
assign MEM[3015] = input_vector[376] << 0;
assign MEM[3016] = -(input_vector[377] << 7);
assign MEM[3017] = input_vector[377] << 6;
assign MEM[3018] = input_vector[377] << 5;
assign MEM[3019] = input_vector[377] << 4;
assign MEM[3020] = input_vector[377] << 3;
assign MEM[3021] = input_vector[377] << 2;
assign MEM[3022] = input_vector[377] << 1;
assign MEM[3023] = input_vector[377] << 0;
assign MEM[3024] = -(input_vector[378] << 7);
assign MEM[3025] = input_vector[378] << 6;
assign MEM[3026] = input_vector[378] << 5;
assign MEM[3027] = input_vector[378] << 4;
assign MEM[3028] = input_vector[378] << 3;
assign MEM[3029] = input_vector[378] << 2;
assign MEM[3030] = input_vector[378] << 1;
assign MEM[3031] = input_vector[378] << 0;
assign MEM[3032] = -(input_vector[379] << 7);
assign MEM[3033] = input_vector[379] << 6;
assign MEM[3034] = input_vector[379] << 5;
assign MEM[3035] = input_vector[379] << 4;
assign MEM[3036] = input_vector[379] << 3;
assign MEM[3037] = input_vector[379] << 2;
assign MEM[3038] = input_vector[379] << 1;
assign MEM[3039] = input_vector[379] << 0;
assign MEM[3040] = -(input_vector[380] << 7);
assign MEM[3041] = input_vector[380] << 6;
assign MEM[3042] = input_vector[380] << 5;
assign MEM[3043] = input_vector[380] << 4;
assign MEM[3044] = input_vector[380] << 3;
assign MEM[3045] = input_vector[380] << 2;
assign MEM[3046] = input_vector[380] << 1;
assign MEM[3047] = input_vector[380] << 0;
assign MEM[3048] = -(input_vector[381] << 7);
assign MEM[3049] = input_vector[381] << 6;
assign MEM[3050] = input_vector[381] << 5;
assign MEM[3051] = input_vector[381] << 4;
assign MEM[3052] = input_vector[381] << 3;
assign MEM[3053] = input_vector[381] << 2;
assign MEM[3054] = input_vector[381] << 1;
assign MEM[3055] = input_vector[381] << 0;
assign MEM[3056] = -(input_vector[382] << 7);
assign MEM[3057] = input_vector[382] << 6;
assign MEM[3058] = input_vector[382] << 5;
assign MEM[3059] = input_vector[382] << 4;
assign MEM[3060] = input_vector[382] << 3;
assign MEM[3061] = input_vector[382] << 2;
assign MEM[3062] = input_vector[382] << 1;
assign MEM[3063] = input_vector[382] << 0;
assign MEM[3064] = -(input_vector[383] << 7);
assign MEM[3065] = input_vector[383] << 6;
assign MEM[3066] = input_vector[383] << 5;
assign MEM[3067] = input_vector[383] << 4;
assign MEM[3068] = input_vector[383] << 3;
assign MEM[3069] = input_vector[383] << 2;
assign MEM[3070] = input_vector[383] << 1;
assign MEM[3071] = input_vector[383] << 0;
assign MEM[3072] = -(input_vector[384] << 7);
assign MEM[3073] = input_vector[384] << 6;
assign MEM[3074] = input_vector[384] << 5;
assign MEM[3075] = input_vector[384] << 4;
assign MEM[3076] = input_vector[384] << 3;
assign MEM[3077] = input_vector[384] << 2;
assign MEM[3078] = input_vector[384] << 1;
assign MEM[3079] = input_vector[384] << 0;
assign MEM[3080] = -(input_vector[385] << 7);
assign MEM[3081] = input_vector[385] << 6;
assign MEM[3082] = input_vector[385] << 5;
assign MEM[3083] = input_vector[385] << 4;
assign MEM[3084] = input_vector[385] << 3;
assign MEM[3085] = input_vector[385] << 2;
assign MEM[3086] = input_vector[385] << 1;
assign MEM[3087] = input_vector[385] << 0;
assign MEM[3088] = -(input_vector[386] << 7);
assign MEM[3089] = input_vector[386] << 6;
assign MEM[3090] = input_vector[386] << 5;
assign MEM[3091] = input_vector[386] << 4;
assign MEM[3092] = input_vector[386] << 3;
assign MEM[3093] = input_vector[386] << 2;
assign MEM[3094] = input_vector[386] << 1;
assign MEM[3095] = input_vector[386] << 0;
assign MEM[3096] = -(input_vector[387] << 7);
assign MEM[3097] = input_vector[387] << 6;
assign MEM[3098] = input_vector[387] << 5;
assign MEM[3099] = input_vector[387] << 4;
assign MEM[3100] = input_vector[387] << 3;
assign MEM[3101] = input_vector[387] << 2;
assign MEM[3102] = input_vector[387] << 1;
assign MEM[3103] = input_vector[387] << 0;
assign MEM[3104] = -(input_vector[388] << 7);
assign MEM[3105] = input_vector[388] << 6;
assign MEM[3106] = input_vector[388] << 5;
assign MEM[3107] = input_vector[388] << 4;
assign MEM[3108] = input_vector[388] << 3;
assign MEM[3109] = input_vector[388] << 2;
assign MEM[3110] = input_vector[388] << 1;
assign MEM[3111] = input_vector[388] << 0;
assign MEM[3112] = -(input_vector[389] << 7);
assign MEM[3113] = input_vector[389] << 6;
assign MEM[3114] = input_vector[389] << 5;
assign MEM[3115] = input_vector[389] << 4;
assign MEM[3116] = input_vector[389] << 3;
assign MEM[3117] = input_vector[389] << 2;
assign MEM[3118] = input_vector[389] << 1;
assign MEM[3119] = input_vector[389] << 0;
assign MEM[3120] = -(input_vector[390] << 7);
assign MEM[3121] = input_vector[390] << 6;
assign MEM[3122] = input_vector[390] << 5;
assign MEM[3123] = input_vector[390] << 4;
assign MEM[3124] = input_vector[390] << 3;
assign MEM[3125] = input_vector[390] << 2;
assign MEM[3126] = input_vector[390] << 1;
assign MEM[3127] = input_vector[390] << 0;
assign MEM[3128] = -(input_vector[391] << 7);
assign MEM[3129] = input_vector[391] << 6;
assign MEM[3130] = input_vector[391] << 5;
assign MEM[3131] = input_vector[391] << 4;
assign MEM[3132] = input_vector[391] << 3;
assign MEM[3133] = input_vector[391] << 2;
assign MEM[3134] = input_vector[391] << 1;
assign MEM[3135] = input_vector[391] << 0;
assign MEM[3136] = -(input_vector[392] << 7);
assign MEM[3137] = input_vector[392] << 6;
assign MEM[3138] = input_vector[392] << 5;
assign MEM[3139] = input_vector[392] << 4;
assign MEM[3140] = input_vector[392] << 3;
assign MEM[3141] = input_vector[392] << 2;
assign MEM[3142] = input_vector[392] << 1;
assign MEM[3143] = input_vector[392] << 0;
assign MEM[3144] = -(input_vector[393] << 7);
assign MEM[3145] = input_vector[393] << 6;
assign MEM[3146] = input_vector[393] << 5;
assign MEM[3147] = input_vector[393] << 4;
assign MEM[3148] = input_vector[393] << 3;
assign MEM[3149] = input_vector[393] << 2;
assign MEM[3150] = input_vector[393] << 1;
assign MEM[3151] = input_vector[393] << 0;
assign MEM[3152] = -(input_vector[394] << 7);
assign MEM[3153] = input_vector[394] << 6;
assign MEM[3154] = input_vector[394] << 5;
assign MEM[3155] = input_vector[394] << 4;
assign MEM[3156] = input_vector[394] << 3;
assign MEM[3157] = input_vector[394] << 2;
assign MEM[3158] = input_vector[394] << 1;
assign MEM[3159] = input_vector[394] << 0;
assign MEM[3160] = -(input_vector[395] << 7);
assign MEM[3161] = input_vector[395] << 6;
assign MEM[3162] = input_vector[395] << 5;
assign MEM[3163] = input_vector[395] << 4;
assign MEM[3164] = input_vector[395] << 3;
assign MEM[3165] = input_vector[395] << 2;
assign MEM[3166] = input_vector[395] << 1;
assign MEM[3167] = input_vector[395] << 0;
assign MEM[3168] = -(input_vector[396] << 7);
assign MEM[3169] = input_vector[396] << 6;
assign MEM[3170] = input_vector[396] << 5;
assign MEM[3171] = input_vector[396] << 4;
assign MEM[3172] = input_vector[396] << 3;
assign MEM[3173] = input_vector[396] << 2;
assign MEM[3174] = input_vector[396] << 1;
assign MEM[3175] = input_vector[396] << 0;
assign MEM[3176] = -(input_vector[397] << 7);
assign MEM[3177] = input_vector[397] << 6;
assign MEM[3178] = input_vector[397] << 5;
assign MEM[3179] = input_vector[397] << 4;
assign MEM[3180] = input_vector[397] << 3;
assign MEM[3181] = input_vector[397] << 2;
assign MEM[3182] = input_vector[397] << 1;
assign MEM[3183] = input_vector[397] << 0;
assign MEM[3184] = -(input_vector[398] << 7);
assign MEM[3185] = input_vector[398] << 6;
assign MEM[3186] = input_vector[398] << 5;
assign MEM[3187] = input_vector[398] << 4;
assign MEM[3188] = input_vector[398] << 3;
assign MEM[3189] = input_vector[398] << 2;
assign MEM[3190] = input_vector[398] << 1;
assign MEM[3191] = input_vector[398] << 0;
assign MEM[3192] = -(input_vector[399] << 7);
assign MEM[3193] = input_vector[399] << 6;
assign MEM[3194] = input_vector[399] << 5;
assign MEM[3195] = input_vector[399] << 4;
assign MEM[3196] = input_vector[399] << 3;
assign MEM[3197] = input_vector[399] << 2;
assign MEM[3198] = input_vector[399] << 1;
assign MEM[3199] = input_vector[399] << 0;
assign MEM[3200] = -(input_vector[400] << 7);
assign MEM[3201] = input_vector[400] << 6;
assign MEM[3202] = input_vector[400] << 5;
assign MEM[3203] = input_vector[400] << 4;
assign MEM[3204] = input_vector[400] << 3;
assign MEM[3205] = input_vector[400] << 2;
assign MEM[3206] = input_vector[400] << 1;
assign MEM[3207] = input_vector[400] << 0;
assign MEM[3208] = -(input_vector[401] << 7);
assign MEM[3209] = input_vector[401] << 6;
assign MEM[3210] = input_vector[401] << 5;
assign MEM[3211] = input_vector[401] << 4;
assign MEM[3212] = input_vector[401] << 3;
assign MEM[3213] = input_vector[401] << 2;
assign MEM[3214] = input_vector[401] << 1;
assign MEM[3215] = input_vector[401] << 0;
assign MEM[3216] = -(input_vector[402] << 7);
assign MEM[3217] = input_vector[402] << 6;
assign MEM[3218] = input_vector[402] << 5;
assign MEM[3219] = input_vector[402] << 4;
assign MEM[3220] = input_vector[402] << 3;
assign MEM[3221] = input_vector[402] << 2;
assign MEM[3222] = input_vector[402] << 1;
assign MEM[3223] = input_vector[402] << 0;
assign MEM[3224] = -(input_vector[403] << 7);
assign MEM[3225] = input_vector[403] << 6;
assign MEM[3226] = input_vector[403] << 5;
assign MEM[3227] = input_vector[403] << 4;
assign MEM[3228] = input_vector[403] << 3;
assign MEM[3229] = input_vector[403] << 2;
assign MEM[3230] = input_vector[403] << 1;
assign MEM[3231] = input_vector[403] << 0;
assign MEM[3232] = -(input_vector[404] << 7);
assign MEM[3233] = input_vector[404] << 6;
assign MEM[3234] = input_vector[404] << 5;
assign MEM[3235] = input_vector[404] << 4;
assign MEM[3236] = input_vector[404] << 3;
assign MEM[3237] = input_vector[404] << 2;
assign MEM[3238] = input_vector[404] << 1;
assign MEM[3239] = input_vector[404] << 0;
assign MEM[3240] = -(input_vector[405] << 7);
assign MEM[3241] = input_vector[405] << 6;
assign MEM[3242] = input_vector[405] << 5;
assign MEM[3243] = input_vector[405] << 4;
assign MEM[3244] = input_vector[405] << 3;
assign MEM[3245] = input_vector[405] << 2;
assign MEM[3246] = input_vector[405] << 1;
assign MEM[3247] = input_vector[405] << 0;
assign MEM[3248] = -(input_vector[406] << 7);
assign MEM[3249] = input_vector[406] << 6;
assign MEM[3250] = input_vector[406] << 5;
assign MEM[3251] = input_vector[406] << 4;
assign MEM[3252] = input_vector[406] << 3;
assign MEM[3253] = input_vector[406] << 2;
assign MEM[3254] = input_vector[406] << 1;
assign MEM[3255] = input_vector[406] << 0;
assign MEM[3256] = -(input_vector[407] << 7);
assign MEM[3257] = input_vector[407] << 6;
assign MEM[3258] = input_vector[407] << 5;
assign MEM[3259] = input_vector[407] << 4;
assign MEM[3260] = input_vector[407] << 3;
assign MEM[3261] = input_vector[407] << 2;
assign MEM[3262] = input_vector[407] << 1;
assign MEM[3263] = input_vector[407] << 0;
assign MEM[3264] = -(input_vector[408] << 7);
assign MEM[3265] = input_vector[408] << 6;
assign MEM[3266] = input_vector[408] << 5;
assign MEM[3267] = input_vector[408] << 4;
assign MEM[3268] = input_vector[408] << 3;
assign MEM[3269] = input_vector[408] << 2;
assign MEM[3270] = input_vector[408] << 1;
assign MEM[3271] = input_vector[408] << 0;
assign MEM[3272] = -(input_vector[409] << 7);
assign MEM[3273] = input_vector[409] << 6;
assign MEM[3274] = input_vector[409] << 5;
assign MEM[3275] = input_vector[409] << 4;
assign MEM[3276] = input_vector[409] << 3;
assign MEM[3277] = input_vector[409] << 2;
assign MEM[3278] = input_vector[409] << 1;
assign MEM[3279] = input_vector[409] << 0;
assign MEM[3280] = -(input_vector[410] << 7);
assign MEM[3281] = input_vector[410] << 6;
assign MEM[3282] = input_vector[410] << 5;
assign MEM[3283] = input_vector[410] << 4;
assign MEM[3284] = input_vector[410] << 3;
assign MEM[3285] = input_vector[410] << 2;
assign MEM[3286] = input_vector[410] << 1;
assign MEM[3287] = input_vector[410] << 0;
assign MEM[3288] = -(input_vector[411] << 7);
assign MEM[3289] = input_vector[411] << 6;
assign MEM[3290] = input_vector[411] << 5;
assign MEM[3291] = input_vector[411] << 4;
assign MEM[3292] = input_vector[411] << 3;
assign MEM[3293] = input_vector[411] << 2;
assign MEM[3294] = input_vector[411] << 1;
assign MEM[3295] = input_vector[411] << 0;
assign MEM[3296] = -(input_vector[412] << 7);
assign MEM[3297] = input_vector[412] << 6;
assign MEM[3298] = input_vector[412] << 5;
assign MEM[3299] = input_vector[412] << 4;
assign MEM[3300] = input_vector[412] << 3;
assign MEM[3301] = input_vector[412] << 2;
assign MEM[3302] = input_vector[412] << 1;
assign MEM[3303] = input_vector[412] << 0;
assign MEM[3304] = -(input_vector[413] << 7);
assign MEM[3305] = input_vector[413] << 6;
assign MEM[3306] = input_vector[413] << 5;
assign MEM[3307] = input_vector[413] << 4;
assign MEM[3308] = input_vector[413] << 3;
assign MEM[3309] = input_vector[413] << 2;
assign MEM[3310] = input_vector[413] << 1;
assign MEM[3311] = input_vector[413] << 0;
assign MEM[3312] = -(input_vector[414] << 7);
assign MEM[3313] = input_vector[414] << 6;
assign MEM[3314] = input_vector[414] << 5;
assign MEM[3315] = input_vector[414] << 4;
assign MEM[3316] = input_vector[414] << 3;
assign MEM[3317] = input_vector[414] << 2;
assign MEM[3318] = input_vector[414] << 1;
assign MEM[3319] = input_vector[414] << 0;
assign MEM[3320] = -(input_vector[415] << 7);
assign MEM[3321] = input_vector[415] << 6;
assign MEM[3322] = input_vector[415] << 5;
assign MEM[3323] = input_vector[415] << 4;
assign MEM[3324] = input_vector[415] << 3;
assign MEM[3325] = input_vector[415] << 2;
assign MEM[3326] = input_vector[415] << 1;
assign MEM[3327] = input_vector[415] << 0;
assign MEM[3328] = -(input_vector[416] << 7);
assign MEM[3329] = input_vector[416] << 6;
assign MEM[3330] = input_vector[416] << 5;
assign MEM[3331] = input_vector[416] << 4;
assign MEM[3332] = input_vector[416] << 3;
assign MEM[3333] = input_vector[416] << 2;
assign MEM[3334] = input_vector[416] << 1;
assign MEM[3335] = input_vector[416] << 0;
assign MEM[3336] = -(input_vector[417] << 7);
assign MEM[3337] = input_vector[417] << 6;
assign MEM[3338] = input_vector[417] << 5;
assign MEM[3339] = input_vector[417] << 4;
assign MEM[3340] = input_vector[417] << 3;
assign MEM[3341] = input_vector[417] << 2;
assign MEM[3342] = input_vector[417] << 1;
assign MEM[3343] = input_vector[417] << 0;
assign MEM[3344] = -(input_vector[418] << 7);
assign MEM[3345] = input_vector[418] << 6;
assign MEM[3346] = input_vector[418] << 5;
assign MEM[3347] = input_vector[418] << 4;
assign MEM[3348] = input_vector[418] << 3;
assign MEM[3349] = input_vector[418] << 2;
assign MEM[3350] = input_vector[418] << 1;
assign MEM[3351] = input_vector[418] << 0;
assign MEM[3352] = -(input_vector[419] << 7);
assign MEM[3353] = input_vector[419] << 6;
assign MEM[3354] = input_vector[419] << 5;
assign MEM[3355] = input_vector[419] << 4;
assign MEM[3356] = input_vector[419] << 3;
assign MEM[3357] = input_vector[419] << 2;
assign MEM[3358] = input_vector[419] << 1;
assign MEM[3359] = input_vector[419] << 0;
assign MEM[3360] = -(input_vector[420] << 7);
assign MEM[3361] = input_vector[420] << 6;
assign MEM[3362] = input_vector[420] << 5;
assign MEM[3363] = input_vector[420] << 4;
assign MEM[3364] = input_vector[420] << 3;
assign MEM[3365] = input_vector[420] << 2;
assign MEM[3366] = input_vector[420] << 1;
assign MEM[3367] = input_vector[420] << 0;
assign MEM[3368] = -(input_vector[421] << 7);
assign MEM[3369] = input_vector[421] << 6;
assign MEM[3370] = input_vector[421] << 5;
assign MEM[3371] = input_vector[421] << 4;
assign MEM[3372] = input_vector[421] << 3;
assign MEM[3373] = input_vector[421] << 2;
assign MEM[3374] = input_vector[421] << 1;
assign MEM[3375] = input_vector[421] << 0;
assign MEM[3376] = -(input_vector[422] << 7);
assign MEM[3377] = input_vector[422] << 6;
assign MEM[3378] = input_vector[422] << 5;
assign MEM[3379] = input_vector[422] << 4;
assign MEM[3380] = input_vector[422] << 3;
assign MEM[3381] = input_vector[422] << 2;
assign MEM[3382] = input_vector[422] << 1;
assign MEM[3383] = input_vector[422] << 0;
assign MEM[3384] = -(input_vector[423] << 7);
assign MEM[3385] = input_vector[423] << 6;
assign MEM[3386] = input_vector[423] << 5;
assign MEM[3387] = input_vector[423] << 4;
assign MEM[3388] = input_vector[423] << 3;
assign MEM[3389] = input_vector[423] << 2;
assign MEM[3390] = input_vector[423] << 1;
assign MEM[3391] = input_vector[423] << 0;
assign MEM[3392] = -(input_vector[424] << 7);
assign MEM[3393] = input_vector[424] << 6;
assign MEM[3394] = input_vector[424] << 5;
assign MEM[3395] = input_vector[424] << 4;
assign MEM[3396] = input_vector[424] << 3;
assign MEM[3397] = input_vector[424] << 2;
assign MEM[3398] = input_vector[424] << 1;
assign MEM[3399] = input_vector[424] << 0;
assign MEM[3400] = -(input_vector[425] << 7);
assign MEM[3401] = input_vector[425] << 6;
assign MEM[3402] = input_vector[425] << 5;
assign MEM[3403] = input_vector[425] << 4;
assign MEM[3404] = input_vector[425] << 3;
assign MEM[3405] = input_vector[425] << 2;
assign MEM[3406] = input_vector[425] << 1;
assign MEM[3407] = input_vector[425] << 0;
assign MEM[3408] = -(input_vector[426] << 7);
assign MEM[3409] = input_vector[426] << 6;
assign MEM[3410] = input_vector[426] << 5;
assign MEM[3411] = input_vector[426] << 4;
assign MEM[3412] = input_vector[426] << 3;
assign MEM[3413] = input_vector[426] << 2;
assign MEM[3414] = input_vector[426] << 1;
assign MEM[3415] = input_vector[426] << 0;
assign MEM[3416] = -(input_vector[427] << 7);
assign MEM[3417] = input_vector[427] << 6;
assign MEM[3418] = input_vector[427] << 5;
assign MEM[3419] = input_vector[427] << 4;
assign MEM[3420] = input_vector[427] << 3;
assign MEM[3421] = input_vector[427] << 2;
assign MEM[3422] = input_vector[427] << 1;
assign MEM[3423] = input_vector[427] << 0;
assign MEM[3424] = -(input_vector[428] << 7);
assign MEM[3425] = input_vector[428] << 6;
assign MEM[3426] = input_vector[428] << 5;
assign MEM[3427] = input_vector[428] << 4;
assign MEM[3428] = input_vector[428] << 3;
assign MEM[3429] = input_vector[428] << 2;
assign MEM[3430] = input_vector[428] << 1;
assign MEM[3431] = input_vector[428] << 0;
assign MEM[3432] = -(input_vector[429] << 7);
assign MEM[3433] = input_vector[429] << 6;
assign MEM[3434] = input_vector[429] << 5;
assign MEM[3435] = input_vector[429] << 4;
assign MEM[3436] = input_vector[429] << 3;
assign MEM[3437] = input_vector[429] << 2;
assign MEM[3438] = input_vector[429] << 1;
assign MEM[3439] = input_vector[429] << 0;
assign MEM[3440] = -(input_vector[430] << 7);
assign MEM[3441] = input_vector[430] << 6;
assign MEM[3442] = input_vector[430] << 5;
assign MEM[3443] = input_vector[430] << 4;
assign MEM[3444] = input_vector[430] << 3;
assign MEM[3445] = input_vector[430] << 2;
assign MEM[3446] = input_vector[430] << 1;
assign MEM[3447] = input_vector[430] << 0;
assign MEM[3448] = -(input_vector[431] << 7);
assign MEM[3449] = input_vector[431] << 6;
assign MEM[3450] = input_vector[431] << 5;
assign MEM[3451] = input_vector[431] << 4;
assign MEM[3452] = input_vector[431] << 3;
assign MEM[3453] = input_vector[431] << 2;
assign MEM[3454] = input_vector[431] << 1;
assign MEM[3455] = input_vector[431] << 0;
assign MEM[3456] = -(input_vector[432] << 7);
assign MEM[3457] = input_vector[432] << 6;
assign MEM[3458] = input_vector[432] << 5;
assign MEM[3459] = input_vector[432] << 4;
assign MEM[3460] = input_vector[432] << 3;
assign MEM[3461] = input_vector[432] << 2;
assign MEM[3462] = input_vector[432] << 1;
assign MEM[3463] = input_vector[432] << 0;
assign MEM[3464] = -(input_vector[433] << 7);
assign MEM[3465] = input_vector[433] << 6;
assign MEM[3466] = input_vector[433] << 5;
assign MEM[3467] = input_vector[433] << 4;
assign MEM[3468] = input_vector[433] << 3;
assign MEM[3469] = input_vector[433] << 2;
assign MEM[3470] = input_vector[433] << 1;
assign MEM[3471] = input_vector[433] << 0;
assign MEM[3472] = -(input_vector[434] << 7);
assign MEM[3473] = input_vector[434] << 6;
assign MEM[3474] = input_vector[434] << 5;
assign MEM[3475] = input_vector[434] << 4;
assign MEM[3476] = input_vector[434] << 3;
assign MEM[3477] = input_vector[434] << 2;
assign MEM[3478] = input_vector[434] << 1;
assign MEM[3479] = input_vector[434] << 0;
assign MEM[3480] = -(input_vector[435] << 7);
assign MEM[3481] = input_vector[435] << 6;
assign MEM[3482] = input_vector[435] << 5;
assign MEM[3483] = input_vector[435] << 4;
assign MEM[3484] = input_vector[435] << 3;
assign MEM[3485] = input_vector[435] << 2;
assign MEM[3486] = input_vector[435] << 1;
assign MEM[3487] = input_vector[435] << 0;
assign MEM[3488] = -(input_vector[436] << 7);
assign MEM[3489] = input_vector[436] << 6;
assign MEM[3490] = input_vector[436] << 5;
assign MEM[3491] = input_vector[436] << 4;
assign MEM[3492] = input_vector[436] << 3;
assign MEM[3493] = input_vector[436] << 2;
assign MEM[3494] = input_vector[436] << 1;
assign MEM[3495] = input_vector[436] << 0;
assign MEM[3496] = -(input_vector[437] << 7);
assign MEM[3497] = input_vector[437] << 6;
assign MEM[3498] = input_vector[437] << 5;
assign MEM[3499] = input_vector[437] << 4;
assign MEM[3500] = input_vector[437] << 3;
assign MEM[3501] = input_vector[437] << 2;
assign MEM[3502] = input_vector[437] << 1;
assign MEM[3503] = input_vector[437] << 0;
assign MEM[3504] = -(input_vector[438] << 7);
assign MEM[3505] = input_vector[438] << 6;
assign MEM[3506] = input_vector[438] << 5;
assign MEM[3507] = input_vector[438] << 4;
assign MEM[3508] = input_vector[438] << 3;
assign MEM[3509] = input_vector[438] << 2;
assign MEM[3510] = input_vector[438] << 1;
assign MEM[3511] = input_vector[438] << 0;
assign MEM[3512] = -(input_vector[439] << 7);
assign MEM[3513] = input_vector[439] << 6;
assign MEM[3514] = input_vector[439] << 5;
assign MEM[3515] = input_vector[439] << 4;
assign MEM[3516] = input_vector[439] << 3;
assign MEM[3517] = input_vector[439] << 2;
assign MEM[3518] = input_vector[439] << 1;
assign MEM[3519] = input_vector[439] << 0;
assign MEM[3520] = -(input_vector[440] << 7);
assign MEM[3521] = input_vector[440] << 6;
assign MEM[3522] = input_vector[440] << 5;
assign MEM[3523] = input_vector[440] << 4;
assign MEM[3524] = input_vector[440] << 3;
assign MEM[3525] = input_vector[440] << 2;
assign MEM[3526] = input_vector[440] << 1;
assign MEM[3527] = input_vector[440] << 0;
assign MEM[3528] = -(input_vector[441] << 7);
assign MEM[3529] = input_vector[441] << 6;
assign MEM[3530] = input_vector[441] << 5;
assign MEM[3531] = input_vector[441] << 4;
assign MEM[3532] = input_vector[441] << 3;
assign MEM[3533] = input_vector[441] << 2;
assign MEM[3534] = input_vector[441] << 1;
assign MEM[3535] = input_vector[441] << 0;
assign MEM[3536] = -(input_vector[442] << 7);
assign MEM[3537] = input_vector[442] << 6;
assign MEM[3538] = input_vector[442] << 5;
assign MEM[3539] = input_vector[442] << 4;
assign MEM[3540] = input_vector[442] << 3;
assign MEM[3541] = input_vector[442] << 2;
assign MEM[3542] = input_vector[442] << 1;
assign MEM[3543] = input_vector[442] << 0;
assign MEM[3544] = -(input_vector[443] << 7);
assign MEM[3545] = input_vector[443] << 6;
assign MEM[3546] = input_vector[443] << 5;
assign MEM[3547] = input_vector[443] << 4;
assign MEM[3548] = input_vector[443] << 3;
assign MEM[3549] = input_vector[443] << 2;
assign MEM[3550] = input_vector[443] << 1;
assign MEM[3551] = input_vector[443] << 0;
assign MEM[3552] = -(input_vector[444] << 7);
assign MEM[3553] = input_vector[444] << 6;
assign MEM[3554] = input_vector[444] << 5;
assign MEM[3555] = input_vector[444] << 4;
assign MEM[3556] = input_vector[444] << 3;
assign MEM[3557] = input_vector[444] << 2;
assign MEM[3558] = input_vector[444] << 1;
assign MEM[3559] = input_vector[444] << 0;
assign MEM[3560] = -(input_vector[445] << 7);
assign MEM[3561] = input_vector[445] << 6;
assign MEM[3562] = input_vector[445] << 5;
assign MEM[3563] = input_vector[445] << 4;
assign MEM[3564] = input_vector[445] << 3;
assign MEM[3565] = input_vector[445] << 2;
assign MEM[3566] = input_vector[445] << 1;
assign MEM[3567] = input_vector[445] << 0;
assign MEM[3568] = -(input_vector[446] << 7);
assign MEM[3569] = input_vector[446] << 6;
assign MEM[3570] = input_vector[446] << 5;
assign MEM[3571] = input_vector[446] << 4;
assign MEM[3572] = input_vector[446] << 3;
assign MEM[3573] = input_vector[446] << 2;
assign MEM[3574] = input_vector[446] << 1;
assign MEM[3575] = input_vector[446] << 0;
assign MEM[3576] = -(input_vector[447] << 7);
assign MEM[3577] = input_vector[447] << 6;
assign MEM[3578] = input_vector[447] << 5;
assign MEM[3579] = input_vector[447] << 4;
assign MEM[3580] = input_vector[447] << 3;
assign MEM[3581] = input_vector[447] << 2;
assign MEM[3582] = input_vector[447] << 1;
assign MEM[3583] = input_vector[447] << 0;
assign MEM[3584] = -(input_vector[448] << 7);
assign MEM[3585] = input_vector[448] << 6;
assign MEM[3586] = input_vector[448] << 5;
assign MEM[3587] = input_vector[448] << 4;
assign MEM[3588] = input_vector[448] << 3;
assign MEM[3589] = input_vector[448] << 2;
assign MEM[3590] = input_vector[448] << 1;
assign MEM[3591] = input_vector[448] << 0;
assign MEM[3592] = -(input_vector[449] << 7);
assign MEM[3593] = input_vector[449] << 6;
assign MEM[3594] = input_vector[449] << 5;
assign MEM[3595] = input_vector[449] << 4;
assign MEM[3596] = input_vector[449] << 3;
assign MEM[3597] = input_vector[449] << 2;
assign MEM[3598] = input_vector[449] << 1;
assign MEM[3599] = input_vector[449] << 0;
assign MEM[3600] = -(input_vector[450] << 7);
assign MEM[3601] = input_vector[450] << 6;
assign MEM[3602] = input_vector[450] << 5;
assign MEM[3603] = input_vector[450] << 4;
assign MEM[3604] = input_vector[450] << 3;
assign MEM[3605] = input_vector[450] << 2;
assign MEM[3606] = input_vector[450] << 1;
assign MEM[3607] = input_vector[450] << 0;
assign MEM[3608] = -(input_vector[451] << 7);
assign MEM[3609] = input_vector[451] << 6;
assign MEM[3610] = input_vector[451] << 5;
assign MEM[3611] = input_vector[451] << 4;
assign MEM[3612] = input_vector[451] << 3;
assign MEM[3613] = input_vector[451] << 2;
assign MEM[3614] = input_vector[451] << 1;
assign MEM[3615] = input_vector[451] << 0;
assign MEM[3616] = -(input_vector[452] << 7);
assign MEM[3617] = input_vector[452] << 6;
assign MEM[3618] = input_vector[452] << 5;
assign MEM[3619] = input_vector[452] << 4;
assign MEM[3620] = input_vector[452] << 3;
assign MEM[3621] = input_vector[452] << 2;
assign MEM[3622] = input_vector[452] << 1;
assign MEM[3623] = input_vector[452] << 0;
assign MEM[3624] = -(input_vector[453] << 7);
assign MEM[3625] = input_vector[453] << 6;
assign MEM[3626] = input_vector[453] << 5;
assign MEM[3627] = input_vector[453] << 4;
assign MEM[3628] = input_vector[453] << 3;
assign MEM[3629] = input_vector[453] << 2;
assign MEM[3630] = input_vector[453] << 1;
assign MEM[3631] = input_vector[453] << 0;
assign MEM[3632] = -(input_vector[454] << 7);
assign MEM[3633] = input_vector[454] << 6;
assign MEM[3634] = input_vector[454] << 5;
assign MEM[3635] = input_vector[454] << 4;
assign MEM[3636] = input_vector[454] << 3;
assign MEM[3637] = input_vector[454] << 2;
assign MEM[3638] = input_vector[454] << 1;
assign MEM[3639] = input_vector[454] << 0;
assign MEM[3640] = -(input_vector[455] << 7);
assign MEM[3641] = input_vector[455] << 6;
assign MEM[3642] = input_vector[455] << 5;
assign MEM[3643] = input_vector[455] << 4;
assign MEM[3644] = input_vector[455] << 3;
assign MEM[3645] = input_vector[455] << 2;
assign MEM[3646] = input_vector[455] << 1;
assign MEM[3647] = input_vector[455] << 0;
assign MEM[3648] = -(input_vector[456] << 7);
assign MEM[3649] = input_vector[456] << 6;
assign MEM[3650] = input_vector[456] << 5;
assign MEM[3651] = input_vector[456] << 4;
assign MEM[3652] = input_vector[456] << 3;
assign MEM[3653] = input_vector[456] << 2;
assign MEM[3654] = input_vector[456] << 1;
assign MEM[3655] = input_vector[456] << 0;
assign MEM[3656] = -(input_vector[457] << 7);
assign MEM[3657] = input_vector[457] << 6;
assign MEM[3658] = input_vector[457] << 5;
assign MEM[3659] = input_vector[457] << 4;
assign MEM[3660] = input_vector[457] << 3;
assign MEM[3661] = input_vector[457] << 2;
assign MEM[3662] = input_vector[457] << 1;
assign MEM[3663] = input_vector[457] << 0;
assign MEM[3664] = -(input_vector[458] << 7);
assign MEM[3665] = input_vector[458] << 6;
assign MEM[3666] = input_vector[458] << 5;
assign MEM[3667] = input_vector[458] << 4;
assign MEM[3668] = input_vector[458] << 3;
assign MEM[3669] = input_vector[458] << 2;
assign MEM[3670] = input_vector[458] << 1;
assign MEM[3671] = input_vector[458] << 0;
assign MEM[3672] = -(input_vector[459] << 7);
assign MEM[3673] = input_vector[459] << 6;
assign MEM[3674] = input_vector[459] << 5;
assign MEM[3675] = input_vector[459] << 4;
assign MEM[3676] = input_vector[459] << 3;
assign MEM[3677] = input_vector[459] << 2;
assign MEM[3678] = input_vector[459] << 1;
assign MEM[3679] = input_vector[459] << 0;
assign MEM[3680] = -(input_vector[460] << 7);
assign MEM[3681] = input_vector[460] << 6;
assign MEM[3682] = input_vector[460] << 5;
assign MEM[3683] = input_vector[460] << 4;
assign MEM[3684] = input_vector[460] << 3;
assign MEM[3685] = input_vector[460] << 2;
assign MEM[3686] = input_vector[460] << 1;
assign MEM[3687] = input_vector[460] << 0;
assign MEM[3688] = -(input_vector[461] << 7);
assign MEM[3689] = input_vector[461] << 6;
assign MEM[3690] = input_vector[461] << 5;
assign MEM[3691] = input_vector[461] << 4;
assign MEM[3692] = input_vector[461] << 3;
assign MEM[3693] = input_vector[461] << 2;
assign MEM[3694] = input_vector[461] << 1;
assign MEM[3695] = input_vector[461] << 0;
assign MEM[3696] = -(input_vector[462] << 7);
assign MEM[3697] = input_vector[462] << 6;
assign MEM[3698] = input_vector[462] << 5;
assign MEM[3699] = input_vector[462] << 4;
assign MEM[3700] = input_vector[462] << 3;
assign MEM[3701] = input_vector[462] << 2;
assign MEM[3702] = input_vector[462] << 1;
assign MEM[3703] = input_vector[462] << 0;
assign MEM[3704] = -(input_vector[463] << 7);
assign MEM[3705] = input_vector[463] << 6;
assign MEM[3706] = input_vector[463] << 5;
assign MEM[3707] = input_vector[463] << 4;
assign MEM[3708] = input_vector[463] << 3;
assign MEM[3709] = input_vector[463] << 2;
assign MEM[3710] = input_vector[463] << 1;
assign MEM[3711] = input_vector[463] << 0;
assign MEM[3712] = -(input_vector[464] << 7);
assign MEM[3713] = input_vector[464] << 6;
assign MEM[3714] = input_vector[464] << 5;
assign MEM[3715] = input_vector[464] << 4;
assign MEM[3716] = input_vector[464] << 3;
assign MEM[3717] = input_vector[464] << 2;
assign MEM[3718] = input_vector[464] << 1;
assign MEM[3719] = input_vector[464] << 0;
assign MEM[3720] = -(input_vector[465] << 7);
assign MEM[3721] = input_vector[465] << 6;
assign MEM[3722] = input_vector[465] << 5;
assign MEM[3723] = input_vector[465] << 4;
assign MEM[3724] = input_vector[465] << 3;
assign MEM[3725] = input_vector[465] << 2;
assign MEM[3726] = input_vector[465] << 1;
assign MEM[3727] = input_vector[465] << 0;
assign MEM[3728] = -(input_vector[466] << 7);
assign MEM[3729] = input_vector[466] << 6;
assign MEM[3730] = input_vector[466] << 5;
assign MEM[3731] = input_vector[466] << 4;
assign MEM[3732] = input_vector[466] << 3;
assign MEM[3733] = input_vector[466] << 2;
assign MEM[3734] = input_vector[466] << 1;
assign MEM[3735] = input_vector[466] << 0;
assign MEM[3736] = -(input_vector[467] << 7);
assign MEM[3737] = input_vector[467] << 6;
assign MEM[3738] = input_vector[467] << 5;
assign MEM[3739] = input_vector[467] << 4;
assign MEM[3740] = input_vector[467] << 3;
assign MEM[3741] = input_vector[467] << 2;
assign MEM[3742] = input_vector[467] << 1;
assign MEM[3743] = input_vector[467] << 0;
assign MEM[3744] = -(input_vector[468] << 7);
assign MEM[3745] = input_vector[468] << 6;
assign MEM[3746] = input_vector[468] << 5;
assign MEM[3747] = input_vector[468] << 4;
assign MEM[3748] = input_vector[468] << 3;
assign MEM[3749] = input_vector[468] << 2;
assign MEM[3750] = input_vector[468] << 1;
assign MEM[3751] = input_vector[468] << 0;
assign MEM[3752] = -(input_vector[469] << 7);
assign MEM[3753] = input_vector[469] << 6;
assign MEM[3754] = input_vector[469] << 5;
assign MEM[3755] = input_vector[469] << 4;
assign MEM[3756] = input_vector[469] << 3;
assign MEM[3757] = input_vector[469] << 2;
assign MEM[3758] = input_vector[469] << 1;
assign MEM[3759] = input_vector[469] << 0;
assign MEM[3760] = -(input_vector[470] << 7);
assign MEM[3761] = input_vector[470] << 6;
assign MEM[3762] = input_vector[470] << 5;
assign MEM[3763] = input_vector[470] << 4;
assign MEM[3764] = input_vector[470] << 3;
assign MEM[3765] = input_vector[470] << 2;
assign MEM[3766] = input_vector[470] << 1;
assign MEM[3767] = input_vector[470] << 0;
assign MEM[3768] = -(input_vector[471] << 7);
assign MEM[3769] = input_vector[471] << 6;
assign MEM[3770] = input_vector[471] << 5;
assign MEM[3771] = input_vector[471] << 4;
assign MEM[3772] = input_vector[471] << 3;
assign MEM[3773] = input_vector[471] << 2;
assign MEM[3774] = input_vector[471] << 1;
assign MEM[3775] = input_vector[471] << 0;
assign MEM[3776] = -(input_vector[472] << 7);
assign MEM[3777] = input_vector[472] << 6;
assign MEM[3778] = input_vector[472] << 5;
assign MEM[3779] = input_vector[472] << 4;
assign MEM[3780] = input_vector[472] << 3;
assign MEM[3781] = input_vector[472] << 2;
assign MEM[3782] = input_vector[472] << 1;
assign MEM[3783] = input_vector[472] << 0;
assign MEM[3784] = -(input_vector[473] << 7);
assign MEM[3785] = input_vector[473] << 6;
assign MEM[3786] = input_vector[473] << 5;
assign MEM[3787] = input_vector[473] << 4;
assign MEM[3788] = input_vector[473] << 3;
assign MEM[3789] = input_vector[473] << 2;
assign MEM[3790] = input_vector[473] << 1;
assign MEM[3791] = input_vector[473] << 0;
assign MEM[3792] = -(input_vector[474] << 7);
assign MEM[3793] = input_vector[474] << 6;
assign MEM[3794] = input_vector[474] << 5;
assign MEM[3795] = input_vector[474] << 4;
assign MEM[3796] = input_vector[474] << 3;
assign MEM[3797] = input_vector[474] << 2;
assign MEM[3798] = input_vector[474] << 1;
assign MEM[3799] = input_vector[474] << 0;
assign MEM[3800] = -(input_vector[475] << 7);
assign MEM[3801] = input_vector[475] << 6;
assign MEM[3802] = input_vector[475] << 5;
assign MEM[3803] = input_vector[475] << 4;
assign MEM[3804] = input_vector[475] << 3;
assign MEM[3805] = input_vector[475] << 2;
assign MEM[3806] = input_vector[475] << 1;
assign MEM[3807] = input_vector[475] << 0;
assign MEM[3808] = -(input_vector[476] << 7);
assign MEM[3809] = input_vector[476] << 6;
assign MEM[3810] = input_vector[476] << 5;
assign MEM[3811] = input_vector[476] << 4;
assign MEM[3812] = input_vector[476] << 3;
assign MEM[3813] = input_vector[476] << 2;
assign MEM[3814] = input_vector[476] << 1;
assign MEM[3815] = input_vector[476] << 0;
assign MEM[3816] = -(input_vector[477] << 7);
assign MEM[3817] = input_vector[477] << 6;
assign MEM[3818] = input_vector[477] << 5;
assign MEM[3819] = input_vector[477] << 4;
assign MEM[3820] = input_vector[477] << 3;
assign MEM[3821] = input_vector[477] << 2;
assign MEM[3822] = input_vector[477] << 1;
assign MEM[3823] = input_vector[477] << 0;
assign MEM[3824] = -(input_vector[478] << 7);
assign MEM[3825] = input_vector[478] << 6;
assign MEM[3826] = input_vector[478] << 5;
assign MEM[3827] = input_vector[478] << 4;
assign MEM[3828] = input_vector[478] << 3;
assign MEM[3829] = input_vector[478] << 2;
assign MEM[3830] = input_vector[478] << 1;
assign MEM[3831] = input_vector[478] << 0;
assign MEM[3832] = -(input_vector[479] << 7);
assign MEM[3833] = input_vector[479] << 6;
assign MEM[3834] = input_vector[479] << 5;
assign MEM[3835] = input_vector[479] << 4;
assign MEM[3836] = input_vector[479] << 3;
assign MEM[3837] = input_vector[479] << 2;
assign MEM[3838] = input_vector[479] << 1;
assign MEM[3839] = input_vector[479] << 0;
assign MEM[3840] = -(input_vector[480] << 7);
assign MEM[3841] = input_vector[480] << 6;
assign MEM[3842] = input_vector[480] << 5;
assign MEM[3843] = input_vector[480] << 4;
assign MEM[3844] = input_vector[480] << 3;
assign MEM[3845] = input_vector[480] << 2;
assign MEM[3846] = input_vector[480] << 1;
assign MEM[3847] = input_vector[480] << 0;
assign MEM[3848] = -(input_vector[481] << 7);
assign MEM[3849] = input_vector[481] << 6;
assign MEM[3850] = input_vector[481] << 5;
assign MEM[3851] = input_vector[481] << 4;
assign MEM[3852] = input_vector[481] << 3;
assign MEM[3853] = input_vector[481] << 2;
assign MEM[3854] = input_vector[481] << 1;
assign MEM[3855] = input_vector[481] << 0;
assign MEM[3856] = -(input_vector[482] << 7);
assign MEM[3857] = input_vector[482] << 6;
assign MEM[3858] = input_vector[482] << 5;
assign MEM[3859] = input_vector[482] << 4;
assign MEM[3860] = input_vector[482] << 3;
assign MEM[3861] = input_vector[482] << 2;
assign MEM[3862] = input_vector[482] << 1;
assign MEM[3863] = input_vector[482] << 0;
assign MEM[3864] = -(input_vector[483] << 7);
assign MEM[3865] = input_vector[483] << 6;
assign MEM[3866] = input_vector[483] << 5;
assign MEM[3867] = input_vector[483] << 4;
assign MEM[3868] = input_vector[483] << 3;
assign MEM[3869] = input_vector[483] << 2;
assign MEM[3870] = input_vector[483] << 1;
assign MEM[3871] = input_vector[483] << 0;
assign MEM[3872] = -(input_vector[484] << 7);
assign MEM[3873] = input_vector[484] << 6;
assign MEM[3874] = input_vector[484] << 5;
assign MEM[3875] = input_vector[484] << 4;
assign MEM[3876] = input_vector[484] << 3;
assign MEM[3877] = input_vector[484] << 2;
assign MEM[3878] = input_vector[484] << 1;
assign MEM[3879] = input_vector[484] << 0;
assign MEM[3880] = -(input_vector[485] << 7);
assign MEM[3881] = input_vector[485] << 6;
assign MEM[3882] = input_vector[485] << 5;
assign MEM[3883] = input_vector[485] << 4;
assign MEM[3884] = input_vector[485] << 3;
assign MEM[3885] = input_vector[485] << 2;
assign MEM[3886] = input_vector[485] << 1;
assign MEM[3887] = input_vector[485] << 0;
assign MEM[3888] = -(input_vector[486] << 7);
assign MEM[3889] = input_vector[486] << 6;
assign MEM[3890] = input_vector[486] << 5;
assign MEM[3891] = input_vector[486] << 4;
assign MEM[3892] = input_vector[486] << 3;
assign MEM[3893] = input_vector[486] << 2;
assign MEM[3894] = input_vector[486] << 1;
assign MEM[3895] = input_vector[486] << 0;
assign MEM[3896] = -(input_vector[487] << 7);
assign MEM[3897] = input_vector[487] << 6;
assign MEM[3898] = input_vector[487] << 5;
assign MEM[3899] = input_vector[487] << 4;
assign MEM[3900] = input_vector[487] << 3;
assign MEM[3901] = input_vector[487] << 2;
assign MEM[3902] = input_vector[487] << 1;
assign MEM[3903] = input_vector[487] << 0;
assign MEM[3904] = -(input_vector[488] << 7);
assign MEM[3905] = input_vector[488] << 6;
assign MEM[3906] = input_vector[488] << 5;
assign MEM[3907] = input_vector[488] << 4;
assign MEM[3908] = input_vector[488] << 3;
assign MEM[3909] = input_vector[488] << 2;
assign MEM[3910] = input_vector[488] << 1;
assign MEM[3911] = input_vector[488] << 0;
assign MEM[3912] = -(input_vector[489] << 7);
assign MEM[3913] = input_vector[489] << 6;
assign MEM[3914] = input_vector[489] << 5;
assign MEM[3915] = input_vector[489] << 4;
assign MEM[3916] = input_vector[489] << 3;
assign MEM[3917] = input_vector[489] << 2;
assign MEM[3918] = input_vector[489] << 1;
assign MEM[3919] = input_vector[489] << 0;
assign MEM[3920] = -(input_vector[490] << 7);
assign MEM[3921] = input_vector[490] << 6;
assign MEM[3922] = input_vector[490] << 5;
assign MEM[3923] = input_vector[490] << 4;
assign MEM[3924] = input_vector[490] << 3;
assign MEM[3925] = input_vector[490] << 2;
assign MEM[3926] = input_vector[490] << 1;
assign MEM[3927] = input_vector[490] << 0;
assign MEM[3928] = -(input_vector[491] << 7);
assign MEM[3929] = input_vector[491] << 6;
assign MEM[3930] = input_vector[491] << 5;
assign MEM[3931] = input_vector[491] << 4;
assign MEM[3932] = input_vector[491] << 3;
assign MEM[3933] = input_vector[491] << 2;
assign MEM[3934] = input_vector[491] << 1;
assign MEM[3935] = input_vector[491] << 0;
assign MEM[3936] = -(input_vector[492] << 7);
assign MEM[3937] = input_vector[492] << 6;
assign MEM[3938] = input_vector[492] << 5;
assign MEM[3939] = input_vector[492] << 4;
assign MEM[3940] = input_vector[492] << 3;
assign MEM[3941] = input_vector[492] << 2;
assign MEM[3942] = input_vector[492] << 1;
assign MEM[3943] = input_vector[492] << 0;
assign MEM[3944] = -(input_vector[493] << 7);
assign MEM[3945] = input_vector[493] << 6;
assign MEM[3946] = input_vector[493] << 5;
assign MEM[3947] = input_vector[493] << 4;
assign MEM[3948] = input_vector[493] << 3;
assign MEM[3949] = input_vector[493] << 2;
assign MEM[3950] = input_vector[493] << 1;
assign MEM[3951] = input_vector[493] << 0;
assign MEM[3952] = -(input_vector[494] << 7);
assign MEM[3953] = input_vector[494] << 6;
assign MEM[3954] = input_vector[494] << 5;
assign MEM[3955] = input_vector[494] << 4;
assign MEM[3956] = input_vector[494] << 3;
assign MEM[3957] = input_vector[494] << 2;
assign MEM[3958] = input_vector[494] << 1;
assign MEM[3959] = input_vector[494] << 0;
assign MEM[3960] = -(input_vector[495] << 7);
assign MEM[3961] = input_vector[495] << 6;
assign MEM[3962] = input_vector[495] << 5;
assign MEM[3963] = input_vector[495] << 4;
assign MEM[3964] = input_vector[495] << 3;
assign MEM[3965] = input_vector[495] << 2;
assign MEM[3966] = input_vector[495] << 1;
assign MEM[3967] = input_vector[495] << 0;
assign MEM[3968] = -(input_vector[496] << 7);
assign MEM[3969] = input_vector[496] << 6;
assign MEM[3970] = input_vector[496] << 5;
assign MEM[3971] = input_vector[496] << 4;
assign MEM[3972] = input_vector[496] << 3;
assign MEM[3973] = input_vector[496] << 2;
assign MEM[3974] = input_vector[496] << 1;
assign MEM[3975] = input_vector[496] << 0;
assign MEM[3976] = -(input_vector[497] << 7);
assign MEM[3977] = input_vector[497] << 6;
assign MEM[3978] = input_vector[497] << 5;
assign MEM[3979] = input_vector[497] << 4;
assign MEM[3980] = input_vector[497] << 3;
assign MEM[3981] = input_vector[497] << 2;
assign MEM[3982] = input_vector[497] << 1;
assign MEM[3983] = input_vector[497] << 0;
assign MEM[3984] = -(input_vector[498] << 7);
assign MEM[3985] = input_vector[498] << 6;
assign MEM[3986] = input_vector[498] << 5;
assign MEM[3987] = input_vector[498] << 4;
assign MEM[3988] = input_vector[498] << 3;
assign MEM[3989] = input_vector[498] << 2;
assign MEM[3990] = input_vector[498] << 1;
assign MEM[3991] = input_vector[498] << 0;
assign MEM[3992] = -(input_vector[499] << 7);
assign MEM[3993] = input_vector[499] << 6;
assign MEM[3994] = input_vector[499] << 5;
assign MEM[3995] = input_vector[499] << 4;
assign MEM[3996] = input_vector[499] << 3;
assign MEM[3997] = input_vector[499] << 2;
assign MEM[3998] = input_vector[499] << 1;
assign MEM[3999] = input_vector[499] << 0;
assign MEM[4000] = -(input_vector[500] << 7);
assign MEM[4001] = input_vector[500] << 6;
assign MEM[4002] = input_vector[500] << 5;
assign MEM[4003] = input_vector[500] << 4;
assign MEM[4004] = input_vector[500] << 3;
assign MEM[4005] = input_vector[500] << 2;
assign MEM[4006] = input_vector[500] << 1;
assign MEM[4007] = input_vector[500] << 0;
assign MEM[4008] = -(input_vector[501] << 7);
assign MEM[4009] = input_vector[501] << 6;
assign MEM[4010] = input_vector[501] << 5;
assign MEM[4011] = input_vector[501] << 4;
assign MEM[4012] = input_vector[501] << 3;
assign MEM[4013] = input_vector[501] << 2;
assign MEM[4014] = input_vector[501] << 1;
assign MEM[4015] = input_vector[501] << 0;
assign MEM[4016] = -(input_vector[502] << 7);
assign MEM[4017] = input_vector[502] << 6;
assign MEM[4018] = input_vector[502] << 5;
assign MEM[4019] = input_vector[502] << 4;
assign MEM[4020] = input_vector[502] << 3;
assign MEM[4021] = input_vector[502] << 2;
assign MEM[4022] = input_vector[502] << 1;
assign MEM[4023] = input_vector[502] << 0;
assign MEM[4024] = -(input_vector[503] << 7);
assign MEM[4025] = input_vector[503] << 6;
assign MEM[4026] = input_vector[503] << 5;
assign MEM[4027] = input_vector[503] << 4;
assign MEM[4028] = input_vector[503] << 3;
assign MEM[4029] = input_vector[503] << 2;
assign MEM[4030] = input_vector[503] << 1;
assign MEM[4031] = input_vector[503] << 0;
assign MEM[4032] = -(input_vector[504] << 7);
assign MEM[4033] = input_vector[504] << 6;
assign MEM[4034] = input_vector[504] << 5;
assign MEM[4035] = input_vector[504] << 4;
assign MEM[4036] = input_vector[504] << 3;
assign MEM[4037] = input_vector[504] << 2;
assign MEM[4038] = input_vector[504] << 1;
assign MEM[4039] = input_vector[504] << 0;
assign MEM[4040] = -(input_vector[505] << 7);
assign MEM[4041] = input_vector[505] << 6;
assign MEM[4042] = input_vector[505] << 5;
assign MEM[4043] = input_vector[505] << 4;
assign MEM[4044] = input_vector[505] << 3;
assign MEM[4045] = input_vector[505] << 2;
assign MEM[4046] = input_vector[505] << 1;
assign MEM[4047] = input_vector[505] << 0;
assign MEM[4048] = -(input_vector[506] << 7);
assign MEM[4049] = input_vector[506] << 6;
assign MEM[4050] = input_vector[506] << 5;
assign MEM[4051] = input_vector[506] << 4;
assign MEM[4052] = input_vector[506] << 3;
assign MEM[4053] = input_vector[506] << 2;
assign MEM[4054] = input_vector[506] << 1;
assign MEM[4055] = input_vector[506] << 0;
assign MEM[4056] = -(input_vector[507] << 7);
assign MEM[4057] = input_vector[507] << 6;
assign MEM[4058] = input_vector[507] << 5;
assign MEM[4059] = input_vector[507] << 4;
assign MEM[4060] = input_vector[507] << 3;
assign MEM[4061] = input_vector[507] << 2;
assign MEM[4062] = input_vector[507] << 1;
assign MEM[4063] = input_vector[507] << 0;
assign MEM[4064] = -(input_vector[508] << 7);
assign MEM[4065] = input_vector[508] << 6;
assign MEM[4066] = input_vector[508] << 5;
assign MEM[4067] = input_vector[508] << 4;
assign MEM[4068] = input_vector[508] << 3;
assign MEM[4069] = input_vector[508] << 2;
assign MEM[4070] = input_vector[508] << 1;
assign MEM[4071] = input_vector[508] << 0;
assign MEM[4072] = -(input_vector[509] << 7);
assign MEM[4073] = input_vector[509] << 6;
assign MEM[4074] = input_vector[509] << 5;
assign MEM[4075] = input_vector[509] << 4;
assign MEM[4076] = input_vector[509] << 3;
assign MEM[4077] = input_vector[509] << 2;
assign MEM[4078] = input_vector[509] << 1;
assign MEM[4079] = input_vector[509] << 0;
assign MEM[4080] = -(input_vector[510] << 7);
assign MEM[4081] = input_vector[510] << 6;
assign MEM[4082] = input_vector[510] << 5;
assign MEM[4083] = input_vector[510] << 4;
assign MEM[4084] = input_vector[510] << 3;
assign MEM[4085] = input_vector[510] << 2;
assign MEM[4086] = input_vector[510] << 1;
assign MEM[4087] = input_vector[510] << 0;
assign MEM[4088] = -(input_vector[511] << 7);
assign MEM[4089] = input_vector[511] << 6;
assign MEM[4090] = input_vector[511] << 5;
assign MEM[4091] = input_vector[511] << 4;
assign MEM[4092] = input_vector[511] << 3;
assign MEM[4093] = input_vector[511] << 2;
assign MEM[4094] = input_vector[511] << 1;
assign MEM[4095] = input_vector[511] << 0;
assign MEM[4096] = -(input_vector[512] << 7);
assign MEM[4097] = input_vector[512] << 6;
assign MEM[4098] = input_vector[512] << 5;
assign MEM[4099] = input_vector[512] << 4;
assign MEM[4100] = input_vector[512] << 3;
assign MEM[4101] = input_vector[512] << 2;
assign MEM[4102] = input_vector[512] << 1;
assign MEM[4103] = input_vector[512] << 0;
assign MEM[4104] = -(input_vector[513] << 7);
assign MEM[4105] = input_vector[513] << 6;
assign MEM[4106] = input_vector[513] << 5;
assign MEM[4107] = input_vector[513] << 4;
assign MEM[4108] = input_vector[513] << 3;
assign MEM[4109] = input_vector[513] << 2;
assign MEM[4110] = input_vector[513] << 1;
assign MEM[4111] = input_vector[513] << 0;
assign MEM[4112] = -(input_vector[514] << 7);
assign MEM[4113] = input_vector[514] << 6;
assign MEM[4114] = input_vector[514] << 5;
assign MEM[4115] = input_vector[514] << 4;
assign MEM[4116] = input_vector[514] << 3;
assign MEM[4117] = input_vector[514] << 2;
assign MEM[4118] = input_vector[514] << 1;
assign MEM[4119] = input_vector[514] << 0;
assign MEM[4120] = -(input_vector[515] << 7);
assign MEM[4121] = input_vector[515] << 6;
assign MEM[4122] = input_vector[515] << 5;
assign MEM[4123] = input_vector[515] << 4;
assign MEM[4124] = input_vector[515] << 3;
assign MEM[4125] = input_vector[515] << 2;
assign MEM[4126] = input_vector[515] << 1;
assign MEM[4127] = input_vector[515] << 0;
assign MEM[4128] = -(input_vector[516] << 7);
assign MEM[4129] = input_vector[516] << 6;
assign MEM[4130] = input_vector[516] << 5;
assign MEM[4131] = input_vector[516] << 4;
assign MEM[4132] = input_vector[516] << 3;
assign MEM[4133] = input_vector[516] << 2;
assign MEM[4134] = input_vector[516] << 1;
assign MEM[4135] = input_vector[516] << 0;
assign MEM[4136] = -(input_vector[517] << 7);
assign MEM[4137] = input_vector[517] << 6;
assign MEM[4138] = input_vector[517] << 5;
assign MEM[4139] = input_vector[517] << 4;
assign MEM[4140] = input_vector[517] << 3;
assign MEM[4141] = input_vector[517] << 2;
assign MEM[4142] = input_vector[517] << 1;
assign MEM[4143] = input_vector[517] << 0;
assign MEM[4144] = -(input_vector[518] << 7);
assign MEM[4145] = input_vector[518] << 6;
assign MEM[4146] = input_vector[518] << 5;
assign MEM[4147] = input_vector[518] << 4;
assign MEM[4148] = input_vector[518] << 3;
assign MEM[4149] = input_vector[518] << 2;
assign MEM[4150] = input_vector[518] << 1;
assign MEM[4151] = input_vector[518] << 0;
assign MEM[4152] = -(input_vector[519] << 7);
assign MEM[4153] = input_vector[519] << 6;
assign MEM[4154] = input_vector[519] << 5;
assign MEM[4155] = input_vector[519] << 4;
assign MEM[4156] = input_vector[519] << 3;
assign MEM[4157] = input_vector[519] << 2;
assign MEM[4158] = input_vector[519] << 1;
assign MEM[4159] = input_vector[519] << 0;
assign MEM[4160] = -(input_vector[520] << 7);
assign MEM[4161] = input_vector[520] << 6;
assign MEM[4162] = input_vector[520] << 5;
assign MEM[4163] = input_vector[520] << 4;
assign MEM[4164] = input_vector[520] << 3;
assign MEM[4165] = input_vector[520] << 2;
assign MEM[4166] = input_vector[520] << 1;
assign MEM[4167] = input_vector[520] << 0;
assign MEM[4168] = -(input_vector[521] << 7);
assign MEM[4169] = input_vector[521] << 6;
assign MEM[4170] = input_vector[521] << 5;
assign MEM[4171] = input_vector[521] << 4;
assign MEM[4172] = input_vector[521] << 3;
assign MEM[4173] = input_vector[521] << 2;
assign MEM[4174] = input_vector[521] << 1;
assign MEM[4175] = input_vector[521] << 0;
assign MEM[4176] = -(input_vector[522] << 7);
assign MEM[4177] = input_vector[522] << 6;
assign MEM[4178] = input_vector[522] << 5;
assign MEM[4179] = input_vector[522] << 4;
assign MEM[4180] = input_vector[522] << 3;
assign MEM[4181] = input_vector[522] << 2;
assign MEM[4182] = input_vector[522] << 1;
assign MEM[4183] = input_vector[522] << 0;
assign MEM[4184] = -(input_vector[523] << 7);
assign MEM[4185] = input_vector[523] << 6;
assign MEM[4186] = input_vector[523] << 5;
assign MEM[4187] = input_vector[523] << 4;
assign MEM[4188] = input_vector[523] << 3;
assign MEM[4189] = input_vector[523] << 2;
assign MEM[4190] = input_vector[523] << 1;
assign MEM[4191] = input_vector[523] << 0;
assign MEM[4192] = -(input_vector[524] << 7);
assign MEM[4193] = input_vector[524] << 6;
assign MEM[4194] = input_vector[524] << 5;
assign MEM[4195] = input_vector[524] << 4;
assign MEM[4196] = input_vector[524] << 3;
assign MEM[4197] = input_vector[524] << 2;
assign MEM[4198] = input_vector[524] << 1;
assign MEM[4199] = input_vector[524] << 0;
assign MEM[4200] = -(input_vector[525] << 7);
assign MEM[4201] = input_vector[525] << 6;
assign MEM[4202] = input_vector[525] << 5;
assign MEM[4203] = input_vector[525] << 4;
assign MEM[4204] = input_vector[525] << 3;
assign MEM[4205] = input_vector[525] << 2;
assign MEM[4206] = input_vector[525] << 1;
assign MEM[4207] = input_vector[525] << 0;
assign MEM[4208] = -(input_vector[526] << 7);
assign MEM[4209] = input_vector[526] << 6;
assign MEM[4210] = input_vector[526] << 5;
assign MEM[4211] = input_vector[526] << 4;
assign MEM[4212] = input_vector[526] << 3;
assign MEM[4213] = input_vector[526] << 2;
assign MEM[4214] = input_vector[526] << 1;
assign MEM[4215] = input_vector[526] << 0;
assign MEM[4216] = -(input_vector[527] << 7);
assign MEM[4217] = input_vector[527] << 6;
assign MEM[4218] = input_vector[527] << 5;
assign MEM[4219] = input_vector[527] << 4;
assign MEM[4220] = input_vector[527] << 3;
assign MEM[4221] = input_vector[527] << 2;
assign MEM[4222] = input_vector[527] << 1;
assign MEM[4223] = input_vector[527] << 0;
assign MEM[4224] = -(input_vector[528] << 7);
assign MEM[4225] = input_vector[528] << 6;
assign MEM[4226] = input_vector[528] << 5;
assign MEM[4227] = input_vector[528] << 4;
assign MEM[4228] = input_vector[528] << 3;
assign MEM[4229] = input_vector[528] << 2;
assign MEM[4230] = input_vector[528] << 1;
assign MEM[4231] = input_vector[528] << 0;
assign MEM[4232] = -(input_vector[529] << 7);
assign MEM[4233] = input_vector[529] << 6;
assign MEM[4234] = input_vector[529] << 5;
assign MEM[4235] = input_vector[529] << 4;
assign MEM[4236] = input_vector[529] << 3;
assign MEM[4237] = input_vector[529] << 2;
assign MEM[4238] = input_vector[529] << 1;
assign MEM[4239] = input_vector[529] << 0;
assign MEM[4240] = -(input_vector[530] << 7);
assign MEM[4241] = input_vector[530] << 6;
assign MEM[4242] = input_vector[530] << 5;
assign MEM[4243] = input_vector[530] << 4;
assign MEM[4244] = input_vector[530] << 3;
assign MEM[4245] = input_vector[530] << 2;
assign MEM[4246] = input_vector[530] << 1;
assign MEM[4247] = input_vector[530] << 0;
assign MEM[4248] = -(input_vector[531] << 7);
assign MEM[4249] = input_vector[531] << 6;
assign MEM[4250] = input_vector[531] << 5;
assign MEM[4251] = input_vector[531] << 4;
assign MEM[4252] = input_vector[531] << 3;
assign MEM[4253] = input_vector[531] << 2;
assign MEM[4254] = input_vector[531] << 1;
assign MEM[4255] = input_vector[531] << 0;
assign MEM[4256] = -(input_vector[532] << 7);
assign MEM[4257] = input_vector[532] << 6;
assign MEM[4258] = input_vector[532] << 5;
assign MEM[4259] = input_vector[532] << 4;
assign MEM[4260] = input_vector[532] << 3;
assign MEM[4261] = input_vector[532] << 2;
assign MEM[4262] = input_vector[532] << 1;
assign MEM[4263] = input_vector[532] << 0;
assign MEM[4264] = -(input_vector[533] << 7);
assign MEM[4265] = input_vector[533] << 6;
assign MEM[4266] = input_vector[533] << 5;
assign MEM[4267] = input_vector[533] << 4;
assign MEM[4268] = input_vector[533] << 3;
assign MEM[4269] = input_vector[533] << 2;
assign MEM[4270] = input_vector[533] << 1;
assign MEM[4271] = input_vector[533] << 0;
assign MEM[4272] = -(input_vector[534] << 7);
assign MEM[4273] = input_vector[534] << 6;
assign MEM[4274] = input_vector[534] << 5;
assign MEM[4275] = input_vector[534] << 4;
assign MEM[4276] = input_vector[534] << 3;
assign MEM[4277] = input_vector[534] << 2;
assign MEM[4278] = input_vector[534] << 1;
assign MEM[4279] = input_vector[534] << 0;
assign MEM[4280] = -(input_vector[535] << 7);
assign MEM[4281] = input_vector[535] << 6;
assign MEM[4282] = input_vector[535] << 5;
assign MEM[4283] = input_vector[535] << 4;
assign MEM[4284] = input_vector[535] << 3;
assign MEM[4285] = input_vector[535] << 2;
assign MEM[4286] = input_vector[535] << 1;
assign MEM[4287] = input_vector[535] << 0;
assign MEM[4288] = -(input_vector[536] << 7);
assign MEM[4289] = input_vector[536] << 6;
assign MEM[4290] = input_vector[536] << 5;
assign MEM[4291] = input_vector[536] << 4;
assign MEM[4292] = input_vector[536] << 3;
assign MEM[4293] = input_vector[536] << 2;
assign MEM[4294] = input_vector[536] << 1;
assign MEM[4295] = input_vector[536] << 0;
assign MEM[4296] = -(input_vector[537] << 7);
assign MEM[4297] = input_vector[537] << 6;
assign MEM[4298] = input_vector[537] << 5;
assign MEM[4299] = input_vector[537] << 4;
assign MEM[4300] = input_vector[537] << 3;
assign MEM[4301] = input_vector[537] << 2;
assign MEM[4302] = input_vector[537] << 1;
assign MEM[4303] = input_vector[537] << 0;
assign MEM[4304] = -(input_vector[538] << 7);
assign MEM[4305] = input_vector[538] << 6;
assign MEM[4306] = input_vector[538] << 5;
assign MEM[4307] = input_vector[538] << 4;
assign MEM[4308] = input_vector[538] << 3;
assign MEM[4309] = input_vector[538] << 2;
assign MEM[4310] = input_vector[538] << 1;
assign MEM[4311] = input_vector[538] << 0;
assign MEM[4312] = -(input_vector[539] << 7);
assign MEM[4313] = input_vector[539] << 6;
assign MEM[4314] = input_vector[539] << 5;
assign MEM[4315] = input_vector[539] << 4;
assign MEM[4316] = input_vector[539] << 3;
assign MEM[4317] = input_vector[539] << 2;
assign MEM[4318] = input_vector[539] << 1;
assign MEM[4319] = input_vector[539] << 0;
assign MEM[4320] = -(input_vector[540] << 7);
assign MEM[4321] = input_vector[540] << 6;
assign MEM[4322] = input_vector[540] << 5;
assign MEM[4323] = input_vector[540] << 4;
assign MEM[4324] = input_vector[540] << 3;
assign MEM[4325] = input_vector[540] << 2;
assign MEM[4326] = input_vector[540] << 1;
assign MEM[4327] = input_vector[540] << 0;
assign MEM[4328] = -(input_vector[541] << 7);
assign MEM[4329] = input_vector[541] << 6;
assign MEM[4330] = input_vector[541] << 5;
assign MEM[4331] = input_vector[541] << 4;
assign MEM[4332] = input_vector[541] << 3;
assign MEM[4333] = input_vector[541] << 2;
assign MEM[4334] = input_vector[541] << 1;
assign MEM[4335] = input_vector[541] << 0;
assign MEM[4336] = -(input_vector[542] << 7);
assign MEM[4337] = input_vector[542] << 6;
assign MEM[4338] = input_vector[542] << 5;
assign MEM[4339] = input_vector[542] << 4;
assign MEM[4340] = input_vector[542] << 3;
assign MEM[4341] = input_vector[542] << 2;
assign MEM[4342] = input_vector[542] << 1;
assign MEM[4343] = input_vector[542] << 0;
assign MEM[4344] = -(input_vector[543] << 7);
assign MEM[4345] = input_vector[543] << 6;
assign MEM[4346] = input_vector[543] << 5;
assign MEM[4347] = input_vector[543] << 4;
assign MEM[4348] = input_vector[543] << 3;
assign MEM[4349] = input_vector[543] << 2;
assign MEM[4350] = input_vector[543] << 1;
assign MEM[4351] = input_vector[543] << 0;
assign MEM[4352] = -(input_vector[544] << 7);
assign MEM[4353] = input_vector[544] << 6;
assign MEM[4354] = input_vector[544] << 5;
assign MEM[4355] = input_vector[544] << 4;
assign MEM[4356] = input_vector[544] << 3;
assign MEM[4357] = input_vector[544] << 2;
assign MEM[4358] = input_vector[544] << 1;
assign MEM[4359] = input_vector[544] << 0;
assign MEM[4360] = -(input_vector[545] << 7);
assign MEM[4361] = input_vector[545] << 6;
assign MEM[4362] = input_vector[545] << 5;
assign MEM[4363] = input_vector[545] << 4;
assign MEM[4364] = input_vector[545] << 3;
assign MEM[4365] = input_vector[545] << 2;
assign MEM[4366] = input_vector[545] << 1;
assign MEM[4367] = input_vector[545] << 0;
assign MEM[4368] = -(input_vector[546] << 7);
assign MEM[4369] = input_vector[546] << 6;
assign MEM[4370] = input_vector[546] << 5;
assign MEM[4371] = input_vector[546] << 4;
assign MEM[4372] = input_vector[546] << 3;
assign MEM[4373] = input_vector[546] << 2;
assign MEM[4374] = input_vector[546] << 1;
assign MEM[4375] = input_vector[546] << 0;
assign MEM[4376] = -(input_vector[547] << 7);
assign MEM[4377] = input_vector[547] << 6;
assign MEM[4378] = input_vector[547] << 5;
assign MEM[4379] = input_vector[547] << 4;
assign MEM[4380] = input_vector[547] << 3;
assign MEM[4381] = input_vector[547] << 2;
assign MEM[4382] = input_vector[547] << 1;
assign MEM[4383] = input_vector[547] << 0;
assign MEM[4384] = -(input_vector[548] << 7);
assign MEM[4385] = input_vector[548] << 6;
assign MEM[4386] = input_vector[548] << 5;
assign MEM[4387] = input_vector[548] << 4;
assign MEM[4388] = input_vector[548] << 3;
assign MEM[4389] = input_vector[548] << 2;
assign MEM[4390] = input_vector[548] << 1;
assign MEM[4391] = input_vector[548] << 0;
assign MEM[4392] = -(input_vector[549] << 7);
assign MEM[4393] = input_vector[549] << 6;
assign MEM[4394] = input_vector[549] << 5;
assign MEM[4395] = input_vector[549] << 4;
assign MEM[4396] = input_vector[549] << 3;
assign MEM[4397] = input_vector[549] << 2;
assign MEM[4398] = input_vector[549] << 1;
assign MEM[4399] = input_vector[549] << 0;
assign MEM[4400] = -(input_vector[550] << 7);
assign MEM[4401] = input_vector[550] << 6;
assign MEM[4402] = input_vector[550] << 5;
assign MEM[4403] = input_vector[550] << 4;
assign MEM[4404] = input_vector[550] << 3;
assign MEM[4405] = input_vector[550] << 2;
assign MEM[4406] = input_vector[550] << 1;
assign MEM[4407] = input_vector[550] << 0;
assign MEM[4408] = -(input_vector[551] << 7);
assign MEM[4409] = input_vector[551] << 6;
assign MEM[4410] = input_vector[551] << 5;
assign MEM[4411] = input_vector[551] << 4;
assign MEM[4412] = input_vector[551] << 3;
assign MEM[4413] = input_vector[551] << 2;
assign MEM[4414] = input_vector[551] << 1;
assign MEM[4415] = input_vector[551] << 0;
assign MEM[4416] = -(input_vector[552] << 7);
assign MEM[4417] = input_vector[552] << 6;
assign MEM[4418] = input_vector[552] << 5;
assign MEM[4419] = input_vector[552] << 4;
assign MEM[4420] = input_vector[552] << 3;
assign MEM[4421] = input_vector[552] << 2;
assign MEM[4422] = input_vector[552] << 1;
assign MEM[4423] = input_vector[552] << 0;
assign MEM[4424] = -(input_vector[553] << 7);
assign MEM[4425] = input_vector[553] << 6;
assign MEM[4426] = input_vector[553] << 5;
assign MEM[4427] = input_vector[553] << 4;
assign MEM[4428] = input_vector[553] << 3;
assign MEM[4429] = input_vector[553] << 2;
assign MEM[4430] = input_vector[553] << 1;
assign MEM[4431] = input_vector[553] << 0;
assign MEM[4432] = -(input_vector[554] << 7);
assign MEM[4433] = input_vector[554] << 6;
assign MEM[4434] = input_vector[554] << 5;
assign MEM[4435] = input_vector[554] << 4;
assign MEM[4436] = input_vector[554] << 3;
assign MEM[4437] = input_vector[554] << 2;
assign MEM[4438] = input_vector[554] << 1;
assign MEM[4439] = input_vector[554] << 0;
assign MEM[4440] = -(input_vector[555] << 7);
assign MEM[4441] = input_vector[555] << 6;
assign MEM[4442] = input_vector[555] << 5;
assign MEM[4443] = input_vector[555] << 4;
assign MEM[4444] = input_vector[555] << 3;
assign MEM[4445] = input_vector[555] << 2;
assign MEM[4446] = input_vector[555] << 1;
assign MEM[4447] = input_vector[555] << 0;
assign MEM[4448] = -(input_vector[556] << 7);
assign MEM[4449] = input_vector[556] << 6;
assign MEM[4450] = input_vector[556] << 5;
assign MEM[4451] = input_vector[556] << 4;
assign MEM[4452] = input_vector[556] << 3;
assign MEM[4453] = input_vector[556] << 2;
assign MEM[4454] = input_vector[556] << 1;
assign MEM[4455] = input_vector[556] << 0;
assign MEM[4456] = -(input_vector[557] << 7);
assign MEM[4457] = input_vector[557] << 6;
assign MEM[4458] = input_vector[557] << 5;
assign MEM[4459] = input_vector[557] << 4;
assign MEM[4460] = input_vector[557] << 3;
assign MEM[4461] = input_vector[557] << 2;
assign MEM[4462] = input_vector[557] << 1;
assign MEM[4463] = input_vector[557] << 0;
assign MEM[4464] = -(input_vector[558] << 7);
assign MEM[4465] = input_vector[558] << 6;
assign MEM[4466] = input_vector[558] << 5;
assign MEM[4467] = input_vector[558] << 4;
assign MEM[4468] = input_vector[558] << 3;
assign MEM[4469] = input_vector[558] << 2;
assign MEM[4470] = input_vector[558] << 1;
assign MEM[4471] = input_vector[558] << 0;
assign MEM[4472] = -(input_vector[559] << 7);
assign MEM[4473] = input_vector[559] << 6;
assign MEM[4474] = input_vector[559] << 5;
assign MEM[4475] = input_vector[559] << 4;
assign MEM[4476] = input_vector[559] << 3;
assign MEM[4477] = input_vector[559] << 2;
assign MEM[4478] = input_vector[559] << 1;
assign MEM[4479] = input_vector[559] << 0;
assign MEM[4480] = -(input_vector[560] << 7);
assign MEM[4481] = input_vector[560] << 6;
assign MEM[4482] = input_vector[560] << 5;
assign MEM[4483] = input_vector[560] << 4;
assign MEM[4484] = input_vector[560] << 3;
assign MEM[4485] = input_vector[560] << 2;
assign MEM[4486] = input_vector[560] << 1;
assign MEM[4487] = input_vector[560] << 0;
assign MEM[4488] = -(input_vector[561] << 7);
assign MEM[4489] = input_vector[561] << 6;
assign MEM[4490] = input_vector[561] << 5;
assign MEM[4491] = input_vector[561] << 4;
assign MEM[4492] = input_vector[561] << 3;
assign MEM[4493] = input_vector[561] << 2;
assign MEM[4494] = input_vector[561] << 1;
assign MEM[4495] = input_vector[561] << 0;
assign MEM[4496] = -(input_vector[562] << 7);
assign MEM[4497] = input_vector[562] << 6;
assign MEM[4498] = input_vector[562] << 5;
assign MEM[4499] = input_vector[562] << 4;
assign MEM[4500] = input_vector[562] << 3;
assign MEM[4501] = input_vector[562] << 2;
assign MEM[4502] = input_vector[562] << 1;
assign MEM[4503] = input_vector[562] << 0;
assign MEM[4504] = -(input_vector[563] << 7);
assign MEM[4505] = input_vector[563] << 6;
assign MEM[4506] = input_vector[563] << 5;
assign MEM[4507] = input_vector[563] << 4;
assign MEM[4508] = input_vector[563] << 3;
assign MEM[4509] = input_vector[563] << 2;
assign MEM[4510] = input_vector[563] << 1;
assign MEM[4511] = input_vector[563] << 0;
assign MEM[4512] = -(input_vector[564] << 7);
assign MEM[4513] = input_vector[564] << 6;
assign MEM[4514] = input_vector[564] << 5;
assign MEM[4515] = input_vector[564] << 4;
assign MEM[4516] = input_vector[564] << 3;
assign MEM[4517] = input_vector[564] << 2;
assign MEM[4518] = input_vector[564] << 1;
assign MEM[4519] = input_vector[564] << 0;
assign MEM[4520] = -(input_vector[565] << 7);
assign MEM[4521] = input_vector[565] << 6;
assign MEM[4522] = input_vector[565] << 5;
assign MEM[4523] = input_vector[565] << 4;
assign MEM[4524] = input_vector[565] << 3;
assign MEM[4525] = input_vector[565] << 2;
assign MEM[4526] = input_vector[565] << 1;
assign MEM[4527] = input_vector[565] << 0;
assign MEM[4528] = -(input_vector[566] << 7);
assign MEM[4529] = input_vector[566] << 6;
assign MEM[4530] = input_vector[566] << 5;
assign MEM[4531] = input_vector[566] << 4;
assign MEM[4532] = input_vector[566] << 3;
assign MEM[4533] = input_vector[566] << 2;
assign MEM[4534] = input_vector[566] << 1;
assign MEM[4535] = input_vector[566] << 0;
assign MEM[4536] = -(input_vector[567] << 7);
assign MEM[4537] = input_vector[567] << 6;
assign MEM[4538] = input_vector[567] << 5;
assign MEM[4539] = input_vector[567] << 4;
assign MEM[4540] = input_vector[567] << 3;
assign MEM[4541] = input_vector[567] << 2;
assign MEM[4542] = input_vector[567] << 1;
assign MEM[4543] = input_vector[567] << 0;
assign MEM[4544] = -(input_vector[568] << 7);
assign MEM[4545] = input_vector[568] << 6;
assign MEM[4546] = input_vector[568] << 5;
assign MEM[4547] = input_vector[568] << 4;
assign MEM[4548] = input_vector[568] << 3;
assign MEM[4549] = input_vector[568] << 2;
assign MEM[4550] = input_vector[568] << 1;
assign MEM[4551] = input_vector[568] << 0;
assign MEM[4552] = -(input_vector[569] << 7);
assign MEM[4553] = input_vector[569] << 6;
assign MEM[4554] = input_vector[569] << 5;
assign MEM[4555] = input_vector[569] << 4;
assign MEM[4556] = input_vector[569] << 3;
assign MEM[4557] = input_vector[569] << 2;
assign MEM[4558] = input_vector[569] << 1;
assign MEM[4559] = input_vector[569] << 0;
assign MEM[4560] = -(input_vector[570] << 7);
assign MEM[4561] = input_vector[570] << 6;
assign MEM[4562] = input_vector[570] << 5;
assign MEM[4563] = input_vector[570] << 4;
assign MEM[4564] = input_vector[570] << 3;
assign MEM[4565] = input_vector[570] << 2;
assign MEM[4566] = input_vector[570] << 1;
assign MEM[4567] = input_vector[570] << 0;
assign MEM[4568] = -(input_vector[571] << 7);
assign MEM[4569] = input_vector[571] << 6;
assign MEM[4570] = input_vector[571] << 5;
assign MEM[4571] = input_vector[571] << 4;
assign MEM[4572] = input_vector[571] << 3;
assign MEM[4573] = input_vector[571] << 2;
assign MEM[4574] = input_vector[571] << 1;
assign MEM[4575] = input_vector[571] << 0;
assign MEM[4576] = -(input_vector[572] << 7);
assign MEM[4577] = input_vector[572] << 6;
assign MEM[4578] = input_vector[572] << 5;
assign MEM[4579] = input_vector[572] << 4;
assign MEM[4580] = input_vector[572] << 3;
assign MEM[4581] = input_vector[572] << 2;
assign MEM[4582] = input_vector[572] << 1;
assign MEM[4583] = input_vector[572] << 0;
assign MEM[4584] = -(input_vector[573] << 7);
assign MEM[4585] = input_vector[573] << 6;
assign MEM[4586] = input_vector[573] << 5;
assign MEM[4587] = input_vector[573] << 4;
assign MEM[4588] = input_vector[573] << 3;
assign MEM[4589] = input_vector[573] << 2;
assign MEM[4590] = input_vector[573] << 1;
assign MEM[4591] = input_vector[573] << 0;
assign MEM[4592] = -(input_vector[574] << 7);
assign MEM[4593] = input_vector[574] << 6;
assign MEM[4594] = input_vector[574] << 5;
assign MEM[4595] = input_vector[574] << 4;
assign MEM[4596] = input_vector[574] << 3;
assign MEM[4597] = input_vector[574] << 2;
assign MEM[4598] = input_vector[574] << 1;
assign MEM[4599] = input_vector[574] << 0;
assign MEM[4600] = -(input_vector[575] << 7);
assign MEM[4601] = input_vector[575] << 6;
assign MEM[4602] = input_vector[575] << 5;
assign MEM[4603] = input_vector[575] << 4;
assign MEM[4604] = input_vector[575] << 3;
assign MEM[4605] = input_vector[575] << 2;
assign MEM[4606] = input_vector[575] << 1;
assign MEM[4607] = input_vector[575] << 0;
assign MEM[4608] = -(input_vector[576] << 7);
assign MEM[4609] = input_vector[576] << 6;
assign MEM[4610] = input_vector[576] << 5;
assign MEM[4611] = input_vector[576] << 4;
assign MEM[4612] = input_vector[576] << 3;
assign MEM[4613] = input_vector[576] << 2;
assign MEM[4614] = input_vector[576] << 1;
assign MEM[4615] = input_vector[576] << 0;
assign MEM[4616] = -(input_vector[577] << 7);
assign MEM[4617] = input_vector[577] << 6;
assign MEM[4618] = input_vector[577] << 5;
assign MEM[4619] = input_vector[577] << 4;
assign MEM[4620] = input_vector[577] << 3;
assign MEM[4621] = input_vector[577] << 2;
assign MEM[4622] = input_vector[577] << 1;
assign MEM[4623] = input_vector[577] << 0;
assign MEM[4624] = -(input_vector[578] << 7);
assign MEM[4625] = input_vector[578] << 6;
assign MEM[4626] = input_vector[578] << 5;
assign MEM[4627] = input_vector[578] << 4;
assign MEM[4628] = input_vector[578] << 3;
assign MEM[4629] = input_vector[578] << 2;
assign MEM[4630] = input_vector[578] << 1;
assign MEM[4631] = input_vector[578] << 0;
assign MEM[4632] = -(input_vector[579] << 7);
assign MEM[4633] = input_vector[579] << 6;
assign MEM[4634] = input_vector[579] << 5;
assign MEM[4635] = input_vector[579] << 4;
assign MEM[4636] = input_vector[579] << 3;
assign MEM[4637] = input_vector[579] << 2;
assign MEM[4638] = input_vector[579] << 1;
assign MEM[4639] = input_vector[579] << 0;
assign MEM[4640] = -(input_vector[580] << 7);
assign MEM[4641] = input_vector[580] << 6;
assign MEM[4642] = input_vector[580] << 5;
assign MEM[4643] = input_vector[580] << 4;
assign MEM[4644] = input_vector[580] << 3;
assign MEM[4645] = input_vector[580] << 2;
assign MEM[4646] = input_vector[580] << 1;
assign MEM[4647] = input_vector[580] << 0;
assign MEM[4648] = -(input_vector[581] << 7);
assign MEM[4649] = input_vector[581] << 6;
assign MEM[4650] = input_vector[581] << 5;
assign MEM[4651] = input_vector[581] << 4;
assign MEM[4652] = input_vector[581] << 3;
assign MEM[4653] = input_vector[581] << 2;
assign MEM[4654] = input_vector[581] << 1;
assign MEM[4655] = input_vector[581] << 0;
assign MEM[4656] = -(input_vector[582] << 7);
assign MEM[4657] = input_vector[582] << 6;
assign MEM[4658] = input_vector[582] << 5;
assign MEM[4659] = input_vector[582] << 4;
assign MEM[4660] = input_vector[582] << 3;
assign MEM[4661] = input_vector[582] << 2;
assign MEM[4662] = input_vector[582] << 1;
assign MEM[4663] = input_vector[582] << 0;
assign MEM[4664] = -(input_vector[583] << 7);
assign MEM[4665] = input_vector[583] << 6;
assign MEM[4666] = input_vector[583] << 5;
assign MEM[4667] = input_vector[583] << 4;
assign MEM[4668] = input_vector[583] << 3;
assign MEM[4669] = input_vector[583] << 2;
assign MEM[4670] = input_vector[583] << 1;
assign MEM[4671] = input_vector[583] << 0;
assign MEM[4672] = -(input_vector[584] << 7);
assign MEM[4673] = input_vector[584] << 6;
assign MEM[4674] = input_vector[584] << 5;
assign MEM[4675] = input_vector[584] << 4;
assign MEM[4676] = input_vector[584] << 3;
assign MEM[4677] = input_vector[584] << 2;
assign MEM[4678] = input_vector[584] << 1;
assign MEM[4679] = input_vector[584] << 0;
assign MEM[4680] = -(input_vector[585] << 7);
assign MEM[4681] = input_vector[585] << 6;
assign MEM[4682] = input_vector[585] << 5;
assign MEM[4683] = input_vector[585] << 4;
assign MEM[4684] = input_vector[585] << 3;
assign MEM[4685] = input_vector[585] << 2;
assign MEM[4686] = input_vector[585] << 1;
assign MEM[4687] = input_vector[585] << 0;
assign MEM[4688] = -(input_vector[586] << 7);
assign MEM[4689] = input_vector[586] << 6;
assign MEM[4690] = input_vector[586] << 5;
assign MEM[4691] = input_vector[586] << 4;
assign MEM[4692] = input_vector[586] << 3;
assign MEM[4693] = input_vector[586] << 2;
assign MEM[4694] = input_vector[586] << 1;
assign MEM[4695] = input_vector[586] << 0;
assign MEM[4696] = -(input_vector[587] << 7);
assign MEM[4697] = input_vector[587] << 6;
assign MEM[4698] = input_vector[587] << 5;
assign MEM[4699] = input_vector[587] << 4;
assign MEM[4700] = input_vector[587] << 3;
assign MEM[4701] = input_vector[587] << 2;
assign MEM[4702] = input_vector[587] << 1;
assign MEM[4703] = input_vector[587] << 0;
assign MEM[4704] = -(input_vector[588] << 7);
assign MEM[4705] = input_vector[588] << 6;
assign MEM[4706] = input_vector[588] << 5;
assign MEM[4707] = input_vector[588] << 4;
assign MEM[4708] = input_vector[588] << 3;
assign MEM[4709] = input_vector[588] << 2;
assign MEM[4710] = input_vector[588] << 1;
assign MEM[4711] = input_vector[588] << 0;
assign MEM[4712] = -(input_vector[589] << 7);
assign MEM[4713] = input_vector[589] << 6;
assign MEM[4714] = input_vector[589] << 5;
assign MEM[4715] = input_vector[589] << 4;
assign MEM[4716] = input_vector[589] << 3;
assign MEM[4717] = input_vector[589] << 2;
assign MEM[4718] = input_vector[589] << 1;
assign MEM[4719] = input_vector[589] << 0;
assign MEM[4720] = -(input_vector[590] << 7);
assign MEM[4721] = input_vector[590] << 6;
assign MEM[4722] = input_vector[590] << 5;
assign MEM[4723] = input_vector[590] << 4;
assign MEM[4724] = input_vector[590] << 3;
assign MEM[4725] = input_vector[590] << 2;
assign MEM[4726] = input_vector[590] << 1;
assign MEM[4727] = input_vector[590] << 0;
assign MEM[4728] = -(input_vector[591] << 7);
assign MEM[4729] = input_vector[591] << 6;
assign MEM[4730] = input_vector[591] << 5;
assign MEM[4731] = input_vector[591] << 4;
assign MEM[4732] = input_vector[591] << 3;
assign MEM[4733] = input_vector[591] << 2;
assign MEM[4734] = input_vector[591] << 1;
assign MEM[4735] = input_vector[591] << 0;
assign MEM[4736] = -(input_vector[592] << 7);
assign MEM[4737] = input_vector[592] << 6;
assign MEM[4738] = input_vector[592] << 5;
assign MEM[4739] = input_vector[592] << 4;
assign MEM[4740] = input_vector[592] << 3;
assign MEM[4741] = input_vector[592] << 2;
assign MEM[4742] = input_vector[592] << 1;
assign MEM[4743] = input_vector[592] << 0;
assign MEM[4744] = -(input_vector[593] << 7);
assign MEM[4745] = input_vector[593] << 6;
assign MEM[4746] = input_vector[593] << 5;
assign MEM[4747] = input_vector[593] << 4;
assign MEM[4748] = input_vector[593] << 3;
assign MEM[4749] = input_vector[593] << 2;
assign MEM[4750] = input_vector[593] << 1;
assign MEM[4751] = input_vector[593] << 0;
assign MEM[4752] = -(input_vector[594] << 7);
assign MEM[4753] = input_vector[594] << 6;
assign MEM[4754] = input_vector[594] << 5;
assign MEM[4755] = input_vector[594] << 4;
assign MEM[4756] = input_vector[594] << 3;
assign MEM[4757] = input_vector[594] << 2;
assign MEM[4758] = input_vector[594] << 1;
assign MEM[4759] = input_vector[594] << 0;
assign MEM[4760] = -(input_vector[595] << 7);
assign MEM[4761] = input_vector[595] << 6;
assign MEM[4762] = input_vector[595] << 5;
assign MEM[4763] = input_vector[595] << 4;
assign MEM[4764] = input_vector[595] << 3;
assign MEM[4765] = input_vector[595] << 2;
assign MEM[4766] = input_vector[595] << 1;
assign MEM[4767] = input_vector[595] << 0;
assign MEM[4768] = -(input_vector[596] << 7);
assign MEM[4769] = input_vector[596] << 6;
assign MEM[4770] = input_vector[596] << 5;
assign MEM[4771] = input_vector[596] << 4;
assign MEM[4772] = input_vector[596] << 3;
assign MEM[4773] = input_vector[596] << 2;
assign MEM[4774] = input_vector[596] << 1;
assign MEM[4775] = input_vector[596] << 0;
assign MEM[4776] = -(input_vector[597] << 7);
assign MEM[4777] = input_vector[597] << 6;
assign MEM[4778] = input_vector[597] << 5;
assign MEM[4779] = input_vector[597] << 4;
assign MEM[4780] = input_vector[597] << 3;
assign MEM[4781] = input_vector[597] << 2;
assign MEM[4782] = input_vector[597] << 1;
assign MEM[4783] = input_vector[597] << 0;
assign MEM[4784] = -(input_vector[598] << 7);
assign MEM[4785] = input_vector[598] << 6;
assign MEM[4786] = input_vector[598] << 5;
assign MEM[4787] = input_vector[598] << 4;
assign MEM[4788] = input_vector[598] << 3;
assign MEM[4789] = input_vector[598] << 2;
assign MEM[4790] = input_vector[598] << 1;
assign MEM[4791] = input_vector[598] << 0;
assign MEM[4792] = -(input_vector[599] << 7);
assign MEM[4793] = input_vector[599] << 6;
assign MEM[4794] = input_vector[599] << 5;
assign MEM[4795] = input_vector[599] << 4;
assign MEM[4796] = input_vector[599] << 3;
assign MEM[4797] = input_vector[599] << 2;
assign MEM[4798] = input_vector[599] << 1;
assign MEM[4799] = input_vector[599] << 0;
assign MEM[4800] = -(input_vector[600] << 7);
assign MEM[4801] = input_vector[600] << 6;
assign MEM[4802] = input_vector[600] << 5;
assign MEM[4803] = input_vector[600] << 4;
assign MEM[4804] = input_vector[600] << 3;
assign MEM[4805] = input_vector[600] << 2;
assign MEM[4806] = input_vector[600] << 1;
assign MEM[4807] = input_vector[600] << 0;
assign MEM[4808] = -(input_vector[601] << 7);
assign MEM[4809] = input_vector[601] << 6;
assign MEM[4810] = input_vector[601] << 5;
assign MEM[4811] = input_vector[601] << 4;
assign MEM[4812] = input_vector[601] << 3;
assign MEM[4813] = input_vector[601] << 2;
assign MEM[4814] = input_vector[601] << 1;
assign MEM[4815] = input_vector[601] << 0;
assign MEM[4816] = -(input_vector[602] << 7);
assign MEM[4817] = input_vector[602] << 6;
assign MEM[4818] = input_vector[602] << 5;
assign MEM[4819] = input_vector[602] << 4;
assign MEM[4820] = input_vector[602] << 3;
assign MEM[4821] = input_vector[602] << 2;
assign MEM[4822] = input_vector[602] << 1;
assign MEM[4823] = input_vector[602] << 0;
assign MEM[4824] = -(input_vector[603] << 7);
assign MEM[4825] = input_vector[603] << 6;
assign MEM[4826] = input_vector[603] << 5;
assign MEM[4827] = input_vector[603] << 4;
assign MEM[4828] = input_vector[603] << 3;
assign MEM[4829] = input_vector[603] << 2;
assign MEM[4830] = input_vector[603] << 1;
assign MEM[4831] = input_vector[603] << 0;
assign MEM[4832] = -(input_vector[604] << 7);
assign MEM[4833] = input_vector[604] << 6;
assign MEM[4834] = input_vector[604] << 5;
assign MEM[4835] = input_vector[604] << 4;
assign MEM[4836] = input_vector[604] << 3;
assign MEM[4837] = input_vector[604] << 2;
assign MEM[4838] = input_vector[604] << 1;
assign MEM[4839] = input_vector[604] << 0;
assign MEM[4840] = -(input_vector[605] << 7);
assign MEM[4841] = input_vector[605] << 6;
assign MEM[4842] = input_vector[605] << 5;
assign MEM[4843] = input_vector[605] << 4;
assign MEM[4844] = input_vector[605] << 3;
assign MEM[4845] = input_vector[605] << 2;
assign MEM[4846] = input_vector[605] << 1;
assign MEM[4847] = input_vector[605] << 0;
assign MEM[4848] = -(input_vector[606] << 7);
assign MEM[4849] = input_vector[606] << 6;
assign MEM[4850] = input_vector[606] << 5;
assign MEM[4851] = input_vector[606] << 4;
assign MEM[4852] = input_vector[606] << 3;
assign MEM[4853] = input_vector[606] << 2;
assign MEM[4854] = input_vector[606] << 1;
assign MEM[4855] = input_vector[606] << 0;
assign MEM[4856] = -(input_vector[607] << 7);
assign MEM[4857] = input_vector[607] << 6;
assign MEM[4858] = input_vector[607] << 5;
assign MEM[4859] = input_vector[607] << 4;
assign MEM[4860] = input_vector[607] << 3;
assign MEM[4861] = input_vector[607] << 2;
assign MEM[4862] = input_vector[607] << 1;
assign MEM[4863] = input_vector[607] << 0;
assign MEM[4864] = -(input_vector[608] << 7);
assign MEM[4865] = input_vector[608] << 6;
assign MEM[4866] = input_vector[608] << 5;
assign MEM[4867] = input_vector[608] << 4;
assign MEM[4868] = input_vector[608] << 3;
assign MEM[4869] = input_vector[608] << 2;
assign MEM[4870] = input_vector[608] << 1;
assign MEM[4871] = input_vector[608] << 0;
assign MEM[4872] = -(input_vector[609] << 7);
assign MEM[4873] = input_vector[609] << 6;
assign MEM[4874] = input_vector[609] << 5;
assign MEM[4875] = input_vector[609] << 4;
assign MEM[4876] = input_vector[609] << 3;
assign MEM[4877] = input_vector[609] << 2;
assign MEM[4878] = input_vector[609] << 1;
assign MEM[4879] = input_vector[609] << 0;
assign MEM[4880] = -(input_vector[610] << 7);
assign MEM[4881] = input_vector[610] << 6;
assign MEM[4882] = input_vector[610] << 5;
assign MEM[4883] = input_vector[610] << 4;
assign MEM[4884] = input_vector[610] << 3;
assign MEM[4885] = input_vector[610] << 2;
assign MEM[4886] = input_vector[610] << 1;
assign MEM[4887] = input_vector[610] << 0;
assign MEM[4888] = -(input_vector[611] << 7);
assign MEM[4889] = input_vector[611] << 6;
assign MEM[4890] = input_vector[611] << 5;
assign MEM[4891] = input_vector[611] << 4;
assign MEM[4892] = input_vector[611] << 3;
assign MEM[4893] = input_vector[611] << 2;
assign MEM[4894] = input_vector[611] << 1;
assign MEM[4895] = input_vector[611] << 0;
assign MEM[4896] = -(input_vector[612] << 7);
assign MEM[4897] = input_vector[612] << 6;
assign MEM[4898] = input_vector[612] << 5;
assign MEM[4899] = input_vector[612] << 4;
assign MEM[4900] = input_vector[612] << 3;
assign MEM[4901] = input_vector[612] << 2;
assign MEM[4902] = input_vector[612] << 1;
assign MEM[4903] = input_vector[612] << 0;
assign MEM[4904] = -(input_vector[613] << 7);
assign MEM[4905] = input_vector[613] << 6;
assign MEM[4906] = input_vector[613] << 5;
assign MEM[4907] = input_vector[613] << 4;
assign MEM[4908] = input_vector[613] << 3;
assign MEM[4909] = input_vector[613] << 2;
assign MEM[4910] = input_vector[613] << 1;
assign MEM[4911] = input_vector[613] << 0;
assign MEM[4912] = -(input_vector[614] << 7);
assign MEM[4913] = input_vector[614] << 6;
assign MEM[4914] = input_vector[614] << 5;
assign MEM[4915] = input_vector[614] << 4;
assign MEM[4916] = input_vector[614] << 3;
assign MEM[4917] = input_vector[614] << 2;
assign MEM[4918] = input_vector[614] << 1;
assign MEM[4919] = input_vector[614] << 0;
assign MEM[4920] = -(input_vector[615] << 7);
assign MEM[4921] = input_vector[615] << 6;
assign MEM[4922] = input_vector[615] << 5;
assign MEM[4923] = input_vector[615] << 4;
assign MEM[4924] = input_vector[615] << 3;
assign MEM[4925] = input_vector[615] << 2;
assign MEM[4926] = input_vector[615] << 1;
assign MEM[4927] = input_vector[615] << 0;
assign MEM[4928] = -(input_vector[616] << 7);
assign MEM[4929] = input_vector[616] << 6;
assign MEM[4930] = input_vector[616] << 5;
assign MEM[4931] = input_vector[616] << 4;
assign MEM[4932] = input_vector[616] << 3;
assign MEM[4933] = input_vector[616] << 2;
assign MEM[4934] = input_vector[616] << 1;
assign MEM[4935] = input_vector[616] << 0;
assign MEM[4936] = -(input_vector[617] << 7);
assign MEM[4937] = input_vector[617] << 6;
assign MEM[4938] = input_vector[617] << 5;
assign MEM[4939] = input_vector[617] << 4;
assign MEM[4940] = input_vector[617] << 3;
assign MEM[4941] = input_vector[617] << 2;
assign MEM[4942] = input_vector[617] << 1;
assign MEM[4943] = input_vector[617] << 0;
assign MEM[4944] = -(input_vector[618] << 7);
assign MEM[4945] = input_vector[618] << 6;
assign MEM[4946] = input_vector[618] << 5;
assign MEM[4947] = input_vector[618] << 4;
assign MEM[4948] = input_vector[618] << 3;
assign MEM[4949] = input_vector[618] << 2;
assign MEM[4950] = input_vector[618] << 1;
assign MEM[4951] = input_vector[618] << 0;
assign MEM[4952] = -(input_vector[619] << 7);
assign MEM[4953] = input_vector[619] << 6;
assign MEM[4954] = input_vector[619] << 5;
assign MEM[4955] = input_vector[619] << 4;
assign MEM[4956] = input_vector[619] << 3;
assign MEM[4957] = input_vector[619] << 2;
assign MEM[4958] = input_vector[619] << 1;
assign MEM[4959] = input_vector[619] << 0;
assign MEM[4960] = -(input_vector[620] << 7);
assign MEM[4961] = input_vector[620] << 6;
assign MEM[4962] = input_vector[620] << 5;
assign MEM[4963] = input_vector[620] << 4;
assign MEM[4964] = input_vector[620] << 3;
assign MEM[4965] = input_vector[620] << 2;
assign MEM[4966] = input_vector[620] << 1;
assign MEM[4967] = input_vector[620] << 0;
assign MEM[4968] = -(input_vector[621] << 7);
assign MEM[4969] = input_vector[621] << 6;
assign MEM[4970] = input_vector[621] << 5;
assign MEM[4971] = input_vector[621] << 4;
assign MEM[4972] = input_vector[621] << 3;
assign MEM[4973] = input_vector[621] << 2;
assign MEM[4974] = input_vector[621] << 1;
assign MEM[4975] = input_vector[621] << 0;
assign MEM[4976] = -(input_vector[622] << 7);
assign MEM[4977] = input_vector[622] << 6;
assign MEM[4978] = input_vector[622] << 5;
assign MEM[4979] = input_vector[622] << 4;
assign MEM[4980] = input_vector[622] << 3;
assign MEM[4981] = input_vector[622] << 2;
assign MEM[4982] = input_vector[622] << 1;
assign MEM[4983] = input_vector[622] << 0;
assign MEM[4984] = -(input_vector[623] << 7);
assign MEM[4985] = input_vector[623] << 6;
assign MEM[4986] = input_vector[623] << 5;
assign MEM[4987] = input_vector[623] << 4;
assign MEM[4988] = input_vector[623] << 3;
assign MEM[4989] = input_vector[623] << 2;
assign MEM[4990] = input_vector[623] << 1;
assign MEM[4991] = input_vector[623] << 0;
assign MEM[4992] = -(input_vector[624] << 7);
assign MEM[4993] = input_vector[624] << 6;
assign MEM[4994] = input_vector[624] << 5;
assign MEM[4995] = input_vector[624] << 4;
assign MEM[4996] = input_vector[624] << 3;
assign MEM[4997] = input_vector[624] << 2;
assign MEM[4998] = input_vector[624] << 1;
assign MEM[4999] = input_vector[624] << 0;
assign MEM[5000] = -(input_vector[625] << 7);
assign MEM[5001] = input_vector[625] << 6;
assign MEM[5002] = input_vector[625] << 5;
assign MEM[5003] = input_vector[625] << 4;
assign MEM[5004] = input_vector[625] << 3;
assign MEM[5005] = input_vector[625] << 2;
assign MEM[5006] = input_vector[625] << 1;
assign MEM[5007] = input_vector[625] << 0;
assign MEM[5008] = -(input_vector[626] << 7);
assign MEM[5009] = input_vector[626] << 6;
assign MEM[5010] = input_vector[626] << 5;
assign MEM[5011] = input_vector[626] << 4;
assign MEM[5012] = input_vector[626] << 3;
assign MEM[5013] = input_vector[626] << 2;
assign MEM[5014] = input_vector[626] << 1;
assign MEM[5015] = input_vector[626] << 0;
assign MEM[5016] = -(input_vector[627] << 7);
assign MEM[5017] = input_vector[627] << 6;
assign MEM[5018] = input_vector[627] << 5;
assign MEM[5019] = input_vector[627] << 4;
assign MEM[5020] = input_vector[627] << 3;
assign MEM[5021] = input_vector[627] << 2;
assign MEM[5022] = input_vector[627] << 1;
assign MEM[5023] = input_vector[627] << 0;
assign MEM[5024] = -(input_vector[628] << 7);
assign MEM[5025] = input_vector[628] << 6;
assign MEM[5026] = input_vector[628] << 5;
assign MEM[5027] = input_vector[628] << 4;
assign MEM[5028] = input_vector[628] << 3;
assign MEM[5029] = input_vector[628] << 2;
assign MEM[5030] = input_vector[628] << 1;
assign MEM[5031] = input_vector[628] << 0;
assign MEM[5032] = -(input_vector[629] << 7);
assign MEM[5033] = input_vector[629] << 6;
assign MEM[5034] = input_vector[629] << 5;
assign MEM[5035] = input_vector[629] << 4;
assign MEM[5036] = input_vector[629] << 3;
assign MEM[5037] = input_vector[629] << 2;
assign MEM[5038] = input_vector[629] << 1;
assign MEM[5039] = input_vector[629] << 0;
assign MEM[5040] = -(input_vector[630] << 7);
assign MEM[5041] = input_vector[630] << 6;
assign MEM[5042] = input_vector[630] << 5;
assign MEM[5043] = input_vector[630] << 4;
assign MEM[5044] = input_vector[630] << 3;
assign MEM[5045] = input_vector[630] << 2;
assign MEM[5046] = input_vector[630] << 1;
assign MEM[5047] = input_vector[630] << 0;
assign MEM[5048] = -(input_vector[631] << 7);
assign MEM[5049] = input_vector[631] << 6;
assign MEM[5050] = input_vector[631] << 5;
assign MEM[5051] = input_vector[631] << 4;
assign MEM[5052] = input_vector[631] << 3;
assign MEM[5053] = input_vector[631] << 2;
assign MEM[5054] = input_vector[631] << 1;
assign MEM[5055] = input_vector[631] << 0;
assign MEM[5056] = -(input_vector[632] << 7);
assign MEM[5057] = input_vector[632] << 6;
assign MEM[5058] = input_vector[632] << 5;
assign MEM[5059] = input_vector[632] << 4;
assign MEM[5060] = input_vector[632] << 3;
assign MEM[5061] = input_vector[632] << 2;
assign MEM[5062] = input_vector[632] << 1;
assign MEM[5063] = input_vector[632] << 0;
assign MEM[5064] = -(input_vector[633] << 7);
assign MEM[5065] = input_vector[633] << 6;
assign MEM[5066] = input_vector[633] << 5;
assign MEM[5067] = input_vector[633] << 4;
assign MEM[5068] = input_vector[633] << 3;
assign MEM[5069] = input_vector[633] << 2;
assign MEM[5070] = input_vector[633] << 1;
assign MEM[5071] = input_vector[633] << 0;
assign MEM[5072] = -(input_vector[634] << 7);
assign MEM[5073] = input_vector[634] << 6;
assign MEM[5074] = input_vector[634] << 5;
assign MEM[5075] = input_vector[634] << 4;
assign MEM[5076] = input_vector[634] << 3;
assign MEM[5077] = input_vector[634] << 2;
assign MEM[5078] = input_vector[634] << 1;
assign MEM[5079] = input_vector[634] << 0;
assign MEM[5080] = -(input_vector[635] << 7);
assign MEM[5081] = input_vector[635] << 6;
assign MEM[5082] = input_vector[635] << 5;
assign MEM[5083] = input_vector[635] << 4;
assign MEM[5084] = input_vector[635] << 3;
assign MEM[5085] = input_vector[635] << 2;
assign MEM[5086] = input_vector[635] << 1;
assign MEM[5087] = input_vector[635] << 0;
assign MEM[5088] = -(input_vector[636] << 7);
assign MEM[5089] = input_vector[636] << 6;
assign MEM[5090] = input_vector[636] << 5;
assign MEM[5091] = input_vector[636] << 4;
assign MEM[5092] = input_vector[636] << 3;
assign MEM[5093] = input_vector[636] << 2;
assign MEM[5094] = input_vector[636] << 1;
assign MEM[5095] = input_vector[636] << 0;
assign MEM[5096] = -(input_vector[637] << 7);
assign MEM[5097] = input_vector[637] << 6;
assign MEM[5098] = input_vector[637] << 5;
assign MEM[5099] = input_vector[637] << 4;
assign MEM[5100] = input_vector[637] << 3;
assign MEM[5101] = input_vector[637] << 2;
assign MEM[5102] = input_vector[637] << 1;
assign MEM[5103] = input_vector[637] << 0;
assign MEM[5104] = -(input_vector[638] << 7);
assign MEM[5105] = input_vector[638] << 6;
assign MEM[5106] = input_vector[638] << 5;
assign MEM[5107] = input_vector[638] << 4;
assign MEM[5108] = input_vector[638] << 3;
assign MEM[5109] = input_vector[638] << 2;
assign MEM[5110] = input_vector[638] << 1;
assign MEM[5111] = input_vector[638] << 0;
assign MEM[5112] = -(input_vector[639] << 7);
assign MEM[5113] = input_vector[639] << 6;
assign MEM[5114] = input_vector[639] << 5;
assign MEM[5115] = input_vector[639] << 4;
assign MEM[5116] = input_vector[639] << 3;
assign MEM[5117] = input_vector[639] << 2;
assign MEM[5118] = input_vector[639] << 1;
assign MEM[5119] = input_vector[639] << 0;
assign MEM[5120] = -(input_vector[640] << 7);
assign MEM[5121] = input_vector[640] << 6;
assign MEM[5122] = input_vector[640] << 5;
assign MEM[5123] = input_vector[640] << 4;
assign MEM[5124] = input_vector[640] << 3;
assign MEM[5125] = input_vector[640] << 2;
assign MEM[5126] = input_vector[640] << 1;
assign MEM[5127] = input_vector[640] << 0;
assign MEM[5128] = -(input_vector[641] << 7);
assign MEM[5129] = input_vector[641] << 6;
assign MEM[5130] = input_vector[641] << 5;
assign MEM[5131] = input_vector[641] << 4;
assign MEM[5132] = input_vector[641] << 3;
assign MEM[5133] = input_vector[641] << 2;
assign MEM[5134] = input_vector[641] << 1;
assign MEM[5135] = input_vector[641] << 0;
assign MEM[5136] = -(input_vector[642] << 7);
assign MEM[5137] = input_vector[642] << 6;
assign MEM[5138] = input_vector[642] << 5;
assign MEM[5139] = input_vector[642] << 4;
assign MEM[5140] = input_vector[642] << 3;
assign MEM[5141] = input_vector[642] << 2;
assign MEM[5142] = input_vector[642] << 1;
assign MEM[5143] = input_vector[642] << 0;
assign MEM[5144] = -(input_vector[643] << 7);
assign MEM[5145] = input_vector[643] << 6;
assign MEM[5146] = input_vector[643] << 5;
assign MEM[5147] = input_vector[643] << 4;
assign MEM[5148] = input_vector[643] << 3;
assign MEM[5149] = input_vector[643] << 2;
assign MEM[5150] = input_vector[643] << 1;
assign MEM[5151] = input_vector[643] << 0;
assign MEM[5152] = -(input_vector[644] << 7);
assign MEM[5153] = input_vector[644] << 6;
assign MEM[5154] = input_vector[644] << 5;
assign MEM[5155] = input_vector[644] << 4;
assign MEM[5156] = input_vector[644] << 3;
assign MEM[5157] = input_vector[644] << 2;
assign MEM[5158] = input_vector[644] << 1;
assign MEM[5159] = input_vector[644] << 0;
assign MEM[5160] = -(input_vector[645] << 7);
assign MEM[5161] = input_vector[645] << 6;
assign MEM[5162] = input_vector[645] << 5;
assign MEM[5163] = input_vector[645] << 4;
assign MEM[5164] = input_vector[645] << 3;
assign MEM[5165] = input_vector[645] << 2;
assign MEM[5166] = input_vector[645] << 1;
assign MEM[5167] = input_vector[645] << 0;
assign MEM[5168] = -(input_vector[646] << 7);
assign MEM[5169] = input_vector[646] << 6;
assign MEM[5170] = input_vector[646] << 5;
assign MEM[5171] = input_vector[646] << 4;
assign MEM[5172] = input_vector[646] << 3;
assign MEM[5173] = input_vector[646] << 2;
assign MEM[5174] = input_vector[646] << 1;
assign MEM[5175] = input_vector[646] << 0;
assign MEM[5176] = -(input_vector[647] << 7);
assign MEM[5177] = input_vector[647] << 6;
assign MEM[5178] = input_vector[647] << 5;
assign MEM[5179] = input_vector[647] << 4;
assign MEM[5180] = input_vector[647] << 3;
assign MEM[5181] = input_vector[647] << 2;
assign MEM[5182] = input_vector[647] << 1;
assign MEM[5183] = input_vector[647] << 0;
assign MEM[5184] = -(input_vector[648] << 7);
assign MEM[5185] = input_vector[648] << 6;
assign MEM[5186] = input_vector[648] << 5;
assign MEM[5187] = input_vector[648] << 4;
assign MEM[5188] = input_vector[648] << 3;
assign MEM[5189] = input_vector[648] << 2;
assign MEM[5190] = input_vector[648] << 1;
assign MEM[5191] = input_vector[648] << 0;
assign MEM[5192] = -(input_vector[649] << 7);
assign MEM[5193] = input_vector[649] << 6;
assign MEM[5194] = input_vector[649] << 5;
assign MEM[5195] = input_vector[649] << 4;
assign MEM[5196] = input_vector[649] << 3;
assign MEM[5197] = input_vector[649] << 2;
assign MEM[5198] = input_vector[649] << 1;
assign MEM[5199] = input_vector[649] << 0;
assign MEM[5200] = -(input_vector[650] << 7);
assign MEM[5201] = input_vector[650] << 6;
assign MEM[5202] = input_vector[650] << 5;
assign MEM[5203] = input_vector[650] << 4;
assign MEM[5204] = input_vector[650] << 3;
assign MEM[5205] = input_vector[650] << 2;
assign MEM[5206] = input_vector[650] << 1;
assign MEM[5207] = input_vector[650] << 0;
assign MEM[5208] = -(input_vector[651] << 7);
assign MEM[5209] = input_vector[651] << 6;
assign MEM[5210] = input_vector[651] << 5;
assign MEM[5211] = input_vector[651] << 4;
assign MEM[5212] = input_vector[651] << 3;
assign MEM[5213] = input_vector[651] << 2;
assign MEM[5214] = input_vector[651] << 1;
assign MEM[5215] = input_vector[651] << 0;
assign MEM[5216] = -(input_vector[652] << 7);
assign MEM[5217] = input_vector[652] << 6;
assign MEM[5218] = input_vector[652] << 5;
assign MEM[5219] = input_vector[652] << 4;
assign MEM[5220] = input_vector[652] << 3;
assign MEM[5221] = input_vector[652] << 2;
assign MEM[5222] = input_vector[652] << 1;
assign MEM[5223] = input_vector[652] << 0;
assign MEM[5224] = -(input_vector[653] << 7);
assign MEM[5225] = input_vector[653] << 6;
assign MEM[5226] = input_vector[653] << 5;
assign MEM[5227] = input_vector[653] << 4;
assign MEM[5228] = input_vector[653] << 3;
assign MEM[5229] = input_vector[653] << 2;
assign MEM[5230] = input_vector[653] << 1;
assign MEM[5231] = input_vector[653] << 0;
assign MEM[5232] = -(input_vector[654] << 7);
assign MEM[5233] = input_vector[654] << 6;
assign MEM[5234] = input_vector[654] << 5;
assign MEM[5235] = input_vector[654] << 4;
assign MEM[5236] = input_vector[654] << 3;
assign MEM[5237] = input_vector[654] << 2;
assign MEM[5238] = input_vector[654] << 1;
assign MEM[5239] = input_vector[654] << 0;
assign MEM[5240] = -(input_vector[655] << 7);
assign MEM[5241] = input_vector[655] << 6;
assign MEM[5242] = input_vector[655] << 5;
assign MEM[5243] = input_vector[655] << 4;
assign MEM[5244] = input_vector[655] << 3;
assign MEM[5245] = input_vector[655] << 2;
assign MEM[5246] = input_vector[655] << 1;
assign MEM[5247] = input_vector[655] << 0;
assign MEM[5248] = -(input_vector[656] << 7);
assign MEM[5249] = input_vector[656] << 6;
assign MEM[5250] = input_vector[656] << 5;
assign MEM[5251] = input_vector[656] << 4;
assign MEM[5252] = input_vector[656] << 3;
assign MEM[5253] = input_vector[656] << 2;
assign MEM[5254] = input_vector[656] << 1;
assign MEM[5255] = input_vector[656] << 0;
assign MEM[5256] = -(input_vector[657] << 7);
assign MEM[5257] = input_vector[657] << 6;
assign MEM[5258] = input_vector[657] << 5;
assign MEM[5259] = input_vector[657] << 4;
assign MEM[5260] = input_vector[657] << 3;
assign MEM[5261] = input_vector[657] << 2;
assign MEM[5262] = input_vector[657] << 1;
assign MEM[5263] = input_vector[657] << 0;
assign MEM[5264] = -(input_vector[658] << 7);
assign MEM[5265] = input_vector[658] << 6;
assign MEM[5266] = input_vector[658] << 5;
assign MEM[5267] = input_vector[658] << 4;
assign MEM[5268] = input_vector[658] << 3;
assign MEM[5269] = input_vector[658] << 2;
assign MEM[5270] = input_vector[658] << 1;
assign MEM[5271] = input_vector[658] << 0;
assign MEM[5272] = -(input_vector[659] << 7);
assign MEM[5273] = input_vector[659] << 6;
assign MEM[5274] = input_vector[659] << 5;
assign MEM[5275] = input_vector[659] << 4;
assign MEM[5276] = input_vector[659] << 3;
assign MEM[5277] = input_vector[659] << 2;
assign MEM[5278] = input_vector[659] << 1;
assign MEM[5279] = input_vector[659] << 0;
assign MEM[5280] = -(input_vector[660] << 7);
assign MEM[5281] = input_vector[660] << 6;
assign MEM[5282] = input_vector[660] << 5;
assign MEM[5283] = input_vector[660] << 4;
assign MEM[5284] = input_vector[660] << 3;
assign MEM[5285] = input_vector[660] << 2;
assign MEM[5286] = input_vector[660] << 1;
assign MEM[5287] = input_vector[660] << 0;
assign MEM[5288] = -(input_vector[661] << 7);
assign MEM[5289] = input_vector[661] << 6;
assign MEM[5290] = input_vector[661] << 5;
assign MEM[5291] = input_vector[661] << 4;
assign MEM[5292] = input_vector[661] << 3;
assign MEM[5293] = input_vector[661] << 2;
assign MEM[5294] = input_vector[661] << 1;
assign MEM[5295] = input_vector[661] << 0;
assign MEM[5296] = -(input_vector[662] << 7);
assign MEM[5297] = input_vector[662] << 6;
assign MEM[5298] = input_vector[662] << 5;
assign MEM[5299] = input_vector[662] << 4;
assign MEM[5300] = input_vector[662] << 3;
assign MEM[5301] = input_vector[662] << 2;
assign MEM[5302] = input_vector[662] << 1;
assign MEM[5303] = input_vector[662] << 0;
assign MEM[5304] = -(input_vector[663] << 7);
assign MEM[5305] = input_vector[663] << 6;
assign MEM[5306] = input_vector[663] << 5;
assign MEM[5307] = input_vector[663] << 4;
assign MEM[5308] = input_vector[663] << 3;
assign MEM[5309] = input_vector[663] << 2;
assign MEM[5310] = input_vector[663] << 1;
assign MEM[5311] = input_vector[663] << 0;
assign MEM[5312] = -(input_vector[664] << 7);
assign MEM[5313] = input_vector[664] << 6;
assign MEM[5314] = input_vector[664] << 5;
assign MEM[5315] = input_vector[664] << 4;
assign MEM[5316] = input_vector[664] << 3;
assign MEM[5317] = input_vector[664] << 2;
assign MEM[5318] = input_vector[664] << 1;
assign MEM[5319] = input_vector[664] << 0;
assign MEM[5320] = -(input_vector[665] << 7);
assign MEM[5321] = input_vector[665] << 6;
assign MEM[5322] = input_vector[665] << 5;
assign MEM[5323] = input_vector[665] << 4;
assign MEM[5324] = input_vector[665] << 3;
assign MEM[5325] = input_vector[665] << 2;
assign MEM[5326] = input_vector[665] << 1;
assign MEM[5327] = input_vector[665] << 0;
assign MEM[5328] = -(input_vector[666] << 7);
assign MEM[5329] = input_vector[666] << 6;
assign MEM[5330] = input_vector[666] << 5;
assign MEM[5331] = input_vector[666] << 4;
assign MEM[5332] = input_vector[666] << 3;
assign MEM[5333] = input_vector[666] << 2;
assign MEM[5334] = input_vector[666] << 1;
assign MEM[5335] = input_vector[666] << 0;
assign MEM[5336] = -(input_vector[667] << 7);
assign MEM[5337] = input_vector[667] << 6;
assign MEM[5338] = input_vector[667] << 5;
assign MEM[5339] = input_vector[667] << 4;
assign MEM[5340] = input_vector[667] << 3;
assign MEM[5341] = input_vector[667] << 2;
assign MEM[5342] = input_vector[667] << 1;
assign MEM[5343] = input_vector[667] << 0;
assign MEM[5344] = -(input_vector[668] << 7);
assign MEM[5345] = input_vector[668] << 6;
assign MEM[5346] = input_vector[668] << 5;
assign MEM[5347] = input_vector[668] << 4;
assign MEM[5348] = input_vector[668] << 3;
assign MEM[5349] = input_vector[668] << 2;
assign MEM[5350] = input_vector[668] << 1;
assign MEM[5351] = input_vector[668] << 0;
assign MEM[5352] = -(input_vector[669] << 7);
assign MEM[5353] = input_vector[669] << 6;
assign MEM[5354] = input_vector[669] << 5;
assign MEM[5355] = input_vector[669] << 4;
assign MEM[5356] = input_vector[669] << 3;
assign MEM[5357] = input_vector[669] << 2;
assign MEM[5358] = input_vector[669] << 1;
assign MEM[5359] = input_vector[669] << 0;
assign MEM[5360] = -(input_vector[670] << 7);
assign MEM[5361] = input_vector[670] << 6;
assign MEM[5362] = input_vector[670] << 5;
assign MEM[5363] = input_vector[670] << 4;
assign MEM[5364] = input_vector[670] << 3;
assign MEM[5365] = input_vector[670] << 2;
assign MEM[5366] = input_vector[670] << 1;
assign MEM[5367] = input_vector[670] << 0;
assign MEM[5368] = -(input_vector[671] << 7);
assign MEM[5369] = input_vector[671] << 6;
assign MEM[5370] = input_vector[671] << 5;
assign MEM[5371] = input_vector[671] << 4;
assign MEM[5372] = input_vector[671] << 3;
assign MEM[5373] = input_vector[671] << 2;
assign MEM[5374] = input_vector[671] << 1;
assign MEM[5375] = input_vector[671] << 0;
assign MEM[5376] = -(input_vector[672] << 7);
assign MEM[5377] = input_vector[672] << 6;
assign MEM[5378] = input_vector[672] << 5;
assign MEM[5379] = input_vector[672] << 4;
assign MEM[5380] = input_vector[672] << 3;
assign MEM[5381] = input_vector[672] << 2;
assign MEM[5382] = input_vector[672] << 1;
assign MEM[5383] = input_vector[672] << 0;
assign MEM[5384] = -(input_vector[673] << 7);
assign MEM[5385] = input_vector[673] << 6;
assign MEM[5386] = input_vector[673] << 5;
assign MEM[5387] = input_vector[673] << 4;
assign MEM[5388] = input_vector[673] << 3;
assign MEM[5389] = input_vector[673] << 2;
assign MEM[5390] = input_vector[673] << 1;
assign MEM[5391] = input_vector[673] << 0;
assign MEM[5392] = -(input_vector[674] << 7);
assign MEM[5393] = input_vector[674] << 6;
assign MEM[5394] = input_vector[674] << 5;
assign MEM[5395] = input_vector[674] << 4;
assign MEM[5396] = input_vector[674] << 3;
assign MEM[5397] = input_vector[674] << 2;
assign MEM[5398] = input_vector[674] << 1;
assign MEM[5399] = input_vector[674] << 0;
assign MEM[5400] = -(input_vector[675] << 7);
assign MEM[5401] = input_vector[675] << 6;
assign MEM[5402] = input_vector[675] << 5;
assign MEM[5403] = input_vector[675] << 4;
assign MEM[5404] = input_vector[675] << 3;
assign MEM[5405] = input_vector[675] << 2;
assign MEM[5406] = input_vector[675] << 1;
assign MEM[5407] = input_vector[675] << 0;
assign MEM[5408] = -(input_vector[676] << 7);
assign MEM[5409] = input_vector[676] << 6;
assign MEM[5410] = input_vector[676] << 5;
assign MEM[5411] = input_vector[676] << 4;
assign MEM[5412] = input_vector[676] << 3;
assign MEM[5413] = input_vector[676] << 2;
assign MEM[5414] = input_vector[676] << 1;
assign MEM[5415] = input_vector[676] << 0;
assign MEM[5416] = -(input_vector[677] << 7);
assign MEM[5417] = input_vector[677] << 6;
assign MEM[5418] = input_vector[677] << 5;
assign MEM[5419] = input_vector[677] << 4;
assign MEM[5420] = input_vector[677] << 3;
assign MEM[5421] = input_vector[677] << 2;
assign MEM[5422] = input_vector[677] << 1;
assign MEM[5423] = input_vector[677] << 0;
assign MEM[5424] = -(input_vector[678] << 7);
assign MEM[5425] = input_vector[678] << 6;
assign MEM[5426] = input_vector[678] << 5;
assign MEM[5427] = input_vector[678] << 4;
assign MEM[5428] = input_vector[678] << 3;
assign MEM[5429] = input_vector[678] << 2;
assign MEM[5430] = input_vector[678] << 1;
assign MEM[5431] = input_vector[678] << 0;
assign MEM[5432] = -(input_vector[679] << 7);
assign MEM[5433] = input_vector[679] << 6;
assign MEM[5434] = input_vector[679] << 5;
assign MEM[5435] = input_vector[679] << 4;
assign MEM[5436] = input_vector[679] << 3;
assign MEM[5437] = input_vector[679] << 2;
assign MEM[5438] = input_vector[679] << 1;
assign MEM[5439] = input_vector[679] << 0;
assign MEM[5440] = -(input_vector[680] << 7);
assign MEM[5441] = input_vector[680] << 6;
assign MEM[5442] = input_vector[680] << 5;
assign MEM[5443] = input_vector[680] << 4;
assign MEM[5444] = input_vector[680] << 3;
assign MEM[5445] = input_vector[680] << 2;
assign MEM[5446] = input_vector[680] << 1;
assign MEM[5447] = input_vector[680] << 0;
assign MEM[5448] = -(input_vector[681] << 7);
assign MEM[5449] = input_vector[681] << 6;
assign MEM[5450] = input_vector[681] << 5;
assign MEM[5451] = input_vector[681] << 4;
assign MEM[5452] = input_vector[681] << 3;
assign MEM[5453] = input_vector[681] << 2;
assign MEM[5454] = input_vector[681] << 1;
assign MEM[5455] = input_vector[681] << 0;
assign MEM[5456] = -(input_vector[682] << 7);
assign MEM[5457] = input_vector[682] << 6;
assign MEM[5458] = input_vector[682] << 5;
assign MEM[5459] = input_vector[682] << 4;
assign MEM[5460] = input_vector[682] << 3;
assign MEM[5461] = input_vector[682] << 2;
assign MEM[5462] = input_vector[682] << 1;
assign MEM[5463] = input_vector[682] << 0;
assign MEM[5464] = -(input_vector[683] << 7);
assign MEM[5465] = input_vector[683] << 6;
assign MEM[5466] = input_vector[683] << 5;
assign MEM[5467] = input_vector[683] << 4;
assign MEM[5468] = input_vector[683] << 3;
assign MEM[5469] = input_vector[683] << 2;
assign MEM[5470] = input_vector[683] << 1;
assign MEM[5471] = input_vector[683] << 0;
assign MEM[5472] = -(input_vector[684] << 7);
assign MEM[5473] = input_vector[684] << 6;
assign MEM[5474] = input_vector[684] << 5;
assign MEM[5475] = input_vector[684] << 4;
assign MEM[5476] = input_vector[684] << 3;
assign MEM[5477] = input_vector[684] << 2;
assign MEM[5478] = input_vector[684] << 1;
assign MEM[5479] = input_vector[684] << 0;
assign MEM[5480] = -(input_vector[685] << 7);
assign MEM[5481] = input_vector[685] << 6;
assign MEM[5482] = input_vector[685] << 5;
assign MEM[5483] = input_vector[685] << 4;
assign MEM[5484] = input_vector[685] << 3;
assign MEM[5485] = input_vector[685] << 2;
assign MEM[5486] = input_vector[685] << 1;
assign MEM[5487] = input_vector[685] << 0;
assign MEM[5488] = -(input_vector[686] << 7);
assign MEM[5489] = input_vector[686] << 6;
assign MEM[5490] = input_vector[686] << 5;
assign MEM[5491] = input_vector[686] << 4;
assign MEM[5492] = input_vector[686] << 3;
assign MEM[5493] = input_vector[686] << 2;
assign MEM[5494] = input_vector[686] << 1;
assign MEM[5495] = input_vector[686] << 0;
assign MEM[5496] = -(input_vector[687] << 7);
assign MEM[5497] = input_vector[687] << 6;
assign MEM[5498] = input_vector[687] << 5;
assign MEM[5499] = input_vector[687] << 4;
assign MEM[5500] = input_vector[687] << 3;
assign MEM[5501] = input_vector[687] << 2;
assign MEM[5502] = input_vector[687] << 1;
assign MEM[5503] = input_vector[687] << 0;
assign MEM[5504] = -(input_vector[688] << 7);
assign MEM[5505] = input_vector[688] << 6;
assign MEM[5506] = input_vector[688] << 5;
assign MEM[5507] = input_vector[688] << 4;
assign MEM[5508] = input_vector[688] << 3;
assign MEM[5509] = input_vector[688] << 2;
assign MEM[5510] = input_vector[688] << 1;
assign MEM[5511] = input_vector[688] << 0;
assign MEM[5512] = -(input_vector[689] << 7);
assign MEM[5513] = input_vector[689] << 6;
assign MEM[5514] = input_vector[689] << 5;
assign MEM[5515] = input_vector[689] << 4;
assign MEM[5516] = input_vector[689] << 3;
assign MEM[5517] = input_vector[689] << 2;
assign MEM[5518] = input_vector[689] << 1;
assign MEM[5519] = input_vector[689] << 0;
assign MEM[5520] = -(input_vector[690] << 7);
assign MEM[5521] = input_vector[690] << 6;
assign MEM[5522] = input_vector[690] << 5;
assign MEM[5523] = input_vector[690] << 4;
assign MEM[5524] = input_vector[690] << 3;
assign MEM[5525] = input_vector[690] << 2;
assign MEM[5526] = input_vector[690] << 1;
assign MEM[5527] = input_vector[690] << 0;
assign MEM[5528] = -(input_vector[691] << 7);
assign MEM[5529] = input_vector[691] << 6;
assign MEM[5530] = input_vector[691] << 5;
assign MEM[5531] = input_vector[691] << 4;
assign MEM[5532] = input_vector[691] << 3;
assign MEM[5533] = input_vector[691] << 2;
assign MEM[5534] = input_vector[691] << 1;
assign MEM[5535] = input_vector[691] << 0;
assign MEM[5536] = -(input_vector[692] << 7);
assign MEM[5537] = input_vector[692] << 6;
assign MEM[5538] = input_vector[692] << 5;
assign MEM[5539] = input_vector[692] << 4;
assign MEM[5540] = input_vector[692] << 3;
assign MEM[5541] = input_vector[692] << 2;
assign MEM[5542] = input_vector[692] << 1;
assign MEM[5543] = input_vector[692] << 0;
assign MEM[5544] = -(input_vector[693] << 7);
assign MEM[5545] = input_vector[693] << 6;
assign MEM[5546] = input_vector[693] << 5;
assign MEM[5547] = input_vector[693] << 4;
assign MEM[5548] = input_vector[693] << 3;
assign MEM[5549] = input_vector[693] << 2;
assign MEM[5550] = input_vector[693] << 1;
assign MEM[5551] = input_vector[693] << 0;
assign MEM[5552] = -(input_vector[694] << 7);
assign MEM[5553] = input_vector[694] << 6;
assign MEM[5554] = input_vector[694] << 5;
assign MEM[5555] = input_vector[694] << 4;
assign MEM[5556] = input_vector[694] << 3;
assign MEM[5557] = input_vector[694] << 2;
assign MEM[5558] = input_vector[694] << 1;
assign MEM[5559] = input_vector[694] << 0;
assign MEM[5560] = -(input_vector[695] << 7);
assign MEM[5561] = input_vector[695] << 6;
assign MEM[5562] = input_vector[695] << 5;
assign MEM[5563] = input_vector[695] << 4;
assign MEM[5564] = input_vector[695] << 3;
assign MEM[5565] = input_vector[695] << 2;
assign MEM[5566] = input_vector[695] << 1;
assign MEM[5567] = input_vector[695] << 0;
assign MEM[5568] = -(input_vector[696] << 7);
assign MEM[5569] = input_vector[696] << 6;
assign MEM[5570] = input_vector[696] << 5;
assign MEM[5571] = input_vector[696] << 4;
assign MEM[5572] = input_vector[696] << 3;
assign MEM[5573] = input_vector[696] << 2;
assign MEM[5574] = input_vector[696] << 1;
assign MEM[5575] = input_vector[696] << 0;
assign MEM[5576] = -(input_vector[697] << 7);
assign MEM[5577] = input_vector[697] << 6;
assign MEM[5578] = input_vector[697] << 5;
assign MEM[5579] = input_vector[697] << 4;
assign MEM[5580] = input_vector[697] << 3;
assign MEM[5581] = input_vector[697] << 2;
assign MEM[5582] = input_vector[697] << 1;
assign MEM[5583] = input_vector[697] << 0;
assign MEM[5584] = -(input_vector[698] << 7);
assign MEM[5585] = input_vector[698] << 6;
assign MEM[5586] = input_vector[698] << 5;
assign MEM[5587] = input_vector[698] << 4;
assign MEM[5588] = input_vector[698] << 3;
assign MEM[5589] = input_vector[698] << 2;
assign MEM[5590] = input_vector[698] << 1;
assign MEM[5591] = input_vector[698] << 0;
assign MEM[5592] = -(input_vector[699] << 7);
assign MEM[5593] = input_vector[699] << 6;
assign MEM[5594] = input_vector[699] << 5;
assign MEM[5595] = input_vector[699] << 4;
assign MEM[5596] = input_vector[699] << 3;
assign MEM[5597] = input_vector[699] << 2;
assign MEM[5598] = input_vector[699] << 1;
assign MEM[5599] = input_vector[699] << 0;
assign MEM[5600] = -(input_vector[700] << 7);
assign MEM[5601] = input_vector[700] << 6;
assign MEM[5602] = input_vector[700] << 5;
assign MEM[5603] = input_vector[700] << 4;
assign MEM[5604] = input_vector[700] << 3;
assign MEM[5605] = input_vector[700] << 2;
assign MEM[5606] = input_vector[700] << 1;
assign MEM[5607] = input_vector[700] << 0;
assign MEM[5608] = -(input_vector[701] << 7);
assign MEM[5609] = input_vector[701] << 6;
assign MEM[5610] = input_vector[701] << 5;
assign MEM[5611] = input_vector[701] << 4;
assign MEM[5612] = input_vector[701] << 3;
assign MEM[5613] = input_vector[701] << 2;
assign MEM[5614] = input_vector[701] << 1;
assign MEM[5615] = input_vector[701] << 0;
assign MEM[5616] = -(input_vector[702] << 7);
assign MEM[5617] = input_vector[702] << 6;
assign MEM[5618] = input_vector[702] << 5;
assign MEM[5619] = input_vector[702] << 4;
assign MEM[5620] = input_vector[702] << 3;
assign MEM[5621] = input_vector[702] << 2;
assign MEM[5622] = input_vector[702] << 1;
assign MEM[5623] = input_vector[702] << 0;
assign MEM[5624] = -(input_vector[703] << 7);
assign MEM[5625] = input_vector[703] << 6;
assign MEM[5626] = input_vector[703] << 5;
assign MEM[5627] = input_vector[703] << 4;
assign MEM[5628] = input_vector[703] << 3;
assign MEM[5629] = input_vector[703] << 2;
assign MEM[5630] = input_vector[703] << 1;
assign MEM[5631] = input_vector[703] << 0;
assign MEM[5632] = -(input_vector[704] << 7);
assign MEM[5633] = input_vector[704] << 6;
assign MEM[5634] = input_vector[704] << 5;
assign MEM[5635] = input_vector[704] << 4;
assign MEM[5636] = input_vector[704] << 3;
assign MEM[5637] = input_vector[704] << 2;
assign MEM[5638] = input_vector[704] << 1;
assign MEM[5639] = input_vector[704] << 0;
assign MEM[5640] = -(input_vector[705] << 7);
assign MEM[5641] = input_vector[705] << 6;
assign MEM[5642] = input_vector[705] << 5;
assign MEM[5643] = input_vector[705] << 4;
assign MEM[5644] = input_vector[705] << 3;
assign MEM[5645] = input_vector[705] << 2;
assign MEM[5646] = input_vector[705] << 1;
assign MEM[5647] = input_vector[705] << 0;
assign MEM[5648] = -(input_vector[706] << 7);
assign MEM[5649] = input_vector[706] << 6;
assign MEM[5650] = input_vector[706] << 5;
assign MEM[5651] = input_vector[706] << 4;
assign MEM[5652] = input_vector[706] << 3;
assign MEM[5653] = input_vector[706] << 2;
assign MEM[5654] = input_vector[706] << 1;
assign MEM[5655] = input_vector[706] << 0;
assign MEM[5656] = -(input_vector[707] << 7);
assign MEM[5657] = input_vector[707] << 6;
assign MEM[5658] = input_vector[707] << 5;
assign MEM[5659] = input_vector[707] << 4;
assign MEM[5660] = input_vector[707] << 3;
assign MEM[5661] = input_vector[707] << 2;
assign MEM[5662] = input_vector[707] << 1;
assign MEM[5663] = input_vector[707] << 0;
assign MEM[5664] = -(input_vector[708] << 7);
assign MEM[5665] = input_vector[708] << 6;
assign MEM[5666] = input_vector[708] << 5;
assign MEM[5667] = input_vector[708] << 4;
assign MEM[5668] = input_vector[708] << 3;
assign MEM[5669] = input_vector[708] << 2;
assign MEM[5670] = input_vector[708] << 1;
assign MEM[5671] = input_vector[708] << 0;
assign MEM[5672] = -(input_vector[709] << 7);
assign MEM[5673] = input_vector[709] << 6;
assign MEM[5674] = input_vector[709] << 5;
assign MEM[5675] = input_vector[709] << 4;
assign MEM[5676] = input_vector[709] << 3;
assign MEM[5677] = input_vector[709] << 2;
assign MEM[5678] = input_vector[709] << 1;
assign MEM[5679] = input_vector[709] << 0;
assign MEM[5680] = -(input_vector[710] << 7);
assign MEM[5681] = input_vector[710] << 6;
assign MEM[5682] = input_vector[710] << 5;
assign MEM[5683] = input_vector[710] << 4;
assign MEM[5684] = input_vector[710] << 3;
assign MEM[5685] = input_vector[710] << 2;
assign MEM[5686] = input_vector[710] << 1;
assign MEM[5687] = input_vector[710] << 0;
assign MEM[5688] = -(input_vector[711] << 7);
assign MEM[5689] = input_vector[711] << 6;
assign MEM[5690] = input_vector[711] << 5;
assign MEM[5691] = input_vector[711] << 4;
assign MEM[5692] = input_vector[711] << 3;
assign MEM[5693] = input_vector[711] << 2;
assign MEM[5694] = input_vector[711] << 1;
assign MEM[5695] = input_vector[711] << 0;
assign MEM[5696] = -(input_vector[712] << 7);
assign MEM[5697] = input_vector[712] << 6;
assign MEM[5698] = input_vector[712] << 5;
assign MEM[5699] = input_vector[712] << 4;
assign MEM[5700] = input_vector[712] << 3;
assign MEM[5701] = input_vector[712] << 2;
assign MEM[5702] = input_vector[712] << 1;
assign MEM[5703] = input_vector[712] << 0;
assign MEM[5704] = -(input_vector[713] << 7);
assign MEM[5705] = input_vector[713] << 6;
assign MEM[5706] = input_vector[713] << 5;
assign MEM[5707] = input_vector[713] << 4;
assign MEM[5708] = input_vector[713] << 3;
assign MEM[5709] = input_vector[713] << 2;
assign MEM[5710] = input_vector[713] << 1;
assign MEM[5711] = input_vector[713] << 0;
assign MEM[5712] = -(input_vector[714] << 7);
assign MEM[5713] = input_vector[714] << 6;
assign MEM[5714] = input_vector[714] << 5;
assign MEM[5715] = input_vector[714] << 4;
assign MEM[5716] = input_vector[714] << 3;
assign MEM[5717] = input_vector[714] << 2;
assign MEM[5718] = input_vector[714] << 1;
assign MEM[5719] = input_vector[714] << 0;
assign MEM[5720] = -(input_vector[715] << 7);
assign MEM[5721] = input_vector[715] << 6;
assign MEM[5722] = input_vector[715] << 5;
assign MEM[5723] = input_vector[715] << 4;
assign MEM[5724] = input_vector[715] << 3;
assign MEM[5725] = input_vector[715] << 2;
assign MEM[5726] = input_vector[715] << 1;
assign MEM[5727] = input_vector[715] << 0;
assign MEM[5728] = -(input_vector[716] << 7);
assign MEM[5729] = input_vector[716] << 6;
assign MEM[5730] = input_vector[716] << 5;
assign MEM[5731] = input_vector[716] << 4;
assign MEM[5732] = input_vector[716] << 3;
assign MEM[5733] = input_vector[716] << 2;
assign MEM[5734] = input_vector[716] << 1;
assign MEM[5735] = input_vector[716] << 0;
assign MEM[5736] = -(input_vector[717] << 7);
assign MEM[5737] = input_vector[717] << 6;
assign MEM[5738] = input_vector[717] << 5;
assign MEM[5739] = input_vector[717] << 4;
assign MEM[5740] = input_vector[717] << 3;
assign MEM[5741] = input_vector[717] << 2;
assign MEM[5742] = input_vector[717] << 1;
assign MEM[5743] = input_vector[717] << 0;
assign MEM[5744] = -(input_vector[718] << 7);
assign MEM[5745] = input_vector[718] << 6;
assign MEM[5746] = input_vector[718] << 5;
assign MEM[5747] = input_vector[718] << 4;
assign MEM[5748] = input_vector[718] << 3;
assign MEM[5749] = input_vector[718] << 2;
assign MEM[5750] = input_vector[718] << 1;
assign MEM[5751] = input_vector[718] << 0;
assign MEM[5752] = -(input_vector[719] << 7);
assign MEM[5753] = input_vector[719] << 6;
assign MEM[5754] = input_vector[719] << 5;
assign MEM[5755] = input_vector[719] << 4;
assign MEM[5756] = input_vector[719] << 3;
assign MEM[5757] = input_vector[719] << 2;
assign MEM[5758] = input_vector[719] << 1;
assign MEM[5759] = input_vector[719] << 0;
assign MEM[5760] = -(input_vector[720] << 7);
assign MEM[5761] = input_vector[720] << 6;
assign MEM[5762] = input_vector[720] << 5;
assign MEM[5763] = input_vector[720] << 4;
assign MEM[5764] = input_vector[720] << 3;
assign MEM[5765] = input_vector[720] << 2;
assign MEM[5766] = input_vector[720] << 1;
assign MEM[5767] = input_vector[720] << 0;
assign MEM[5768] = -(input_vector[721] << 7);
assign MEM[5769] = input_vector[721] << 6;
assign MEM[5770] = input_vector[721] << 5;
assign MEM[5771] = input_vector[721] << 4;
assign MEM[5772] = input_vector[721] << 3;
assign MEM[5773] = input_vector[721] << 2;
assign MEM[5774] = input_vector[721] << 1;
assign MEM[5775] = input_vector[721] << 0;
assign MEM[5776] = -(input_vector[722] << 7);
assign MEM[5777] = input_vector[722] << 6;
assign MEM[5778] = input_vector[722] << 5;
assign MEM[5779] = input_vector[722] << 4;
assign MEM[5780] = input_vector[722] << 3;
assign MEM[5781] = input_vector[722] << 2;
assign MEM[5782] = input_vector[722] << 1;
assign MEM[5783] = input_vector[722] << 0;
assign MEM[5784] = -(input_vector[723] << 7);
assign MEM[5785] = input_vector[723] << 6;
assign MEM[5786] = input_vector[723] << 5;
assign MEM[5787] = input_vector[723] << 4;
assign MEM[5788] = input_vector[723] << 3;
assign MEM[5789] = input_vector[723] << 2;
assign MEM[5790] = input_vector[723] << 1;
assign MEM[5791] = input_vector[723] << 0;
assign MEM[5792] = -(input_vector[724] << 7);
assign MEM[5793] = input_vector[724] << 6;
assign MEM[5794] = input_vector[724] << 5;
assign MEM[5795] = input_vector[724] << 4;
assign MEM[5796] = input_vector[724] << 3;
assign MEM[5797] = input_vector[724] << 2;
assign MEM[5798] = input_vector[724] << 1;
assign MEM[5799] = input_vector[724] << 0;
assign MEM[5800] = -(input_vector[725] << 7);
assign MEM[5801] = input_vector[725] << 6;
assign MEM[5802] = input_vector[725] << 5;
assign MEM[5803] = input_vector[725] << 4;
assign MEM[5804] = input_vector[725] << 3;
assign MEM[5805] = input_vector[725] << 2;
assign MEM[5806] = input_vector[725] << 1;
assign MEM[5807] = input_vector[725] << 0;
assign MEM[5808] = -(input_vector[726] << 7);
assign MEM[5809] = input_vector[726] << 6;
assign MEM[5810] = input_vector[726] << 5;
assign MEM[5811] = input_vector[726] << 4;
assign MEM[5812] = input_vector[726] << 3;
assign MEM[5813] = input_vector[726] << 2;
assign MEM[5814] = input_vector[726] << 1;
assign MEM[5815] = input_vector[726] << 0;
assign MEM[5816] = -(input_vector[727] << 7);
assign MEM[5817] = input_vector[727] << 6;
assign MEM[5818] = input_vector[727] << 5;
assign MEM[5819] = input_vector[727] << 4;
assign MEM[5820] = input_vector[727] << 3;
assign MEM[5821] = input_vector[727] << 2;
assign MEM[5822] = input_vector[727] << 1;
assign MEM[5823] = input_vector[727] << 0;
assign MEM[5824] = -(input_vector[728] << 7);
assign MEM[5825] = input_vector[728] << 6;
assign MEM[5826] = input_vector[728] << 5;
assign MEM[5827] = input_vector[728] << 4;
assign MEM[5828] = input_vector[728] << 3;
assign MEM[5829] = input_vector[728] << 2;
assign MEM[5830] = input_vector[728] << 1;
assign MEM[5831] = input_vector[728] << 0;
assign MEM[5832] = -(input_vector[729] << 7);
assign MEM[5833] = input_vector[729] << 6;
assign MEM[5834] = input_vector[729] << 5;
assign MEM[5835] = input_vector[729] << 4;
assign MEM[5836] = input_vector[729] << 3;
assign MEM[5837] = input_vector[729] << 2;
assign MEM[5838] = input_vector[729] << 1;
assign MEM[5839] = input_vector[729] << 0;
assign MEM[5840] = -(input_vector[730] << 7);
assign MEM[5841] = input_vector[730] << 6;
assign MEM[5842] = input_vector[730] << 5;
assign MEM[5843] = input_vector[730] << 4;
assign MEM[5844] = input_vector[730] << 3;
assign MEM[5845] = input_vector[730] << 2;
assign MEM[5846] = input_vector[730] << 1;
assign MEM[5847] = input_vector[730] << 0;
assign MEM[5848] = -(input_vector[731] << 7);
assign MEM[5849] = input_vector[731] << 6;
assign MEM[5850] = input_vector[731] << 5;
assign MEM[5851] = input_vector[731] << 4;
assign MEM[5852] = input_vector[731] << 3;
assign MEM[5853] = input_vector[731] << 2;
assign MEM[5854] = input_vector[731] << 1;
assign MEM[5855] = input_vector[731] << 0;
assign MEM[5856] = -(input_vector[732] << 7);
assign MEM[5857] = input_vector[732] << 6;
assign MEM[5858] = input_vector[732] << 5;
assign MEM[5859] = input_vector[732] << 4;
assign MEM[5860] = input_vector[732] << 3;
assign MEM[5861] = input_vector[732] << 2;
assign MEM[5862] = input_vector[732] << 1;
assign MEM[5863] = input_vector[732] << 0;
assign MEM[5864] = -(input_vector[733] << 7);
assign MEM[5865] = input_vector[733] << 6;
assign MEM[5866] = input_vector[733] << 5;
assign MEM[5867] = input_vector[733] << 4;
assign MEM[5868] = input_vector[733] << 3;
assign MEM[5869] = input_vector[733] << 2;
assign MEM[5870] = input_vector[733] << 1;
assign MEM[5871] = input_vector[733] << 0;
assign MEM[5872] = -(input_vector[734] << 7);
assign MEM[5873] = input_vector[734] << 6;
assign MEM[5874] = input_vector[734] << 5;
assign MEM[5875] = input_vector[734] << 4;
assign MEM[5876] = input_vector[734] << 3;
assign MEM[5877] = input_vector[734] << 2;
assign MEM[5878] = input_vector[734] << 1;
assign MEM[5879] = input_vector[734] << 0;
assign MEM[5880] = -(input_vector[735] << 7);
assign MEM[5881] = input_vector[735] << 6;
assign MEM[5882] = input_vector[735] << 5;
assign MEM[5883] = input_vector[735] << 4;
assign MEM[5884] = input_vector[735] << 3;
assign MEM[5885] = input_vector[735] << 2;
assign MEM[5886] = input_vector[735] << 1;
assign MEM[5887] = input_vector[735] << 0;
assign MEM[5888] = -(input_vector[736] << 7);
assign MEM[5889] = input_vector[736] << 6;
assign MEM[5890] = input_vector[736] << 5;
assign MEM[5891] = input_vector[736] << 4;
assign MEM[5892] = input_vector[736] << 3;
assign MEM[5893] = input_vector[736] << 2;
assign MEM[5894] = input_vector[736] << 1;
assign MEM[5895] = input_vector[736] << 0;
assign MEM[5896] = -(input_vector[737] << 7);
assign MEM[5897] = input_vector[737] << 6;
assign MEM[5898] = input_vector[737] << 5;
assign MEM[5899] = input_vector[737] << 4;
assign MEM[5900] = input_vector[737] << 3;
assign MEM[5901] = input_vector[737] << 2;
assign MEM[5902] = input_vector[737] << 1;
assign MEM[5903] = input_vector[737] << 0;
assign MEM[5904] = -(input_vector[738] << 7);
assign MEM[5905] = input_vector[738] << 6;
assign MEM[5906] = input_vector[738] << 5;
assign MEM[5907] = input_vector[738] << 4;
assign MEM[5908] = input_vector[738] << 3;
assign MEM[5909] = input_vector[738] << 2;
assign MEM[5910] = input_vector[738] << 1;
assign MEM[5911] = input_vector[738] << 0;
assign MEM[5912] = -(input_vector[739] << 7);
assign MEM[5913] = input_vector[739] << 6;
assign MEM[5914] = input_vector[739] << 5;
assign MEM[5915] = input_vector[739] << 4;
assign MEM[5916] = input_vector[739] << 3;
assign MEM[5917] = input_vector[739] << 2;
assign MEM[5918] = input_vector[739] << 1;
assign MEM[5919] = input_vector[739] << 0;
assign MEM[5920] = -(input_vector[740] << 7);
assign MEM[5921] = input_vector[740] << 6;
assign MEM[5922] = input_vector[740] << 5;
assign MEM[5923] = input_vector[740] << 4;
assign MEM[5924] = input_vector[740] << 3;
assign MEM[5925] = input_vector[740] << 2;
assign MEM[5926] = input_vector[740] << 1;
assign MEM[5927] = input_vector[740] << 0;
assign MEM[5928] = -(input_vector[741] << 7);
assign MEM[5929] = input_vector[741] << 6;
assign MEM[5930] = input_vector[741] << 5;
assign MEM[5931] = input_vector[741] << 4;
assign MEM[5932] = input_vector[741] << 3;
assign MEM[5933] = input_vector[741] << 2;
assign MEM[5934] = input_vector[741] << 1;
assign MEM[5935] = input_vector[741] << 0;
assign MEM[5936] = -(input_vector[742] << 7);
assign MEM[5937] = input_vector[742] << 6;
assign MEM[5938] = input_vector[742] << 5;
assign MEM[5939] = input_vector[742] << 4;
assign MEM[5940] = input_vector[742] << 3;
assign MEM[5941] = input_vector[742] << 2;
assign MEM[5942] = input_vector[742] << 1;
assign MEM[5943] = input_vector[742] << 0;
assign MEM[5944] = -(input_vector[743] << 7);
assign MEM[5945] = input_vector[743] << 6;
assign MEM[5946] = input_vector[743] << 5;
assign MEM[5947] = input_vector[743] << 4;
assign MEM[5948] = input_vector[743] << 3;
assign MEM[5949] = input_vector[743] << 2;
assign MEM[5950] = input_vector[743] << 1;
assign MEM[5951] = input_vector[743] << 0;
assign MEM[5952] = -(input_vector[744] << 7);
assign MEM[5953] = input_vector[744] << 6;
assign MEM[5954] = input_vector[744] << 5;
assign MEM[5955] = input_vector[744] << 4;
assign MEM[5956] = input_vector[744] << 3;
assign MEM[5957] = input_vector[744] << 2;
assign MEM[5958] = input_vector[744] << 1;
assign MEM[5959] = input_vector[744] << 0;
assign MEM[5960] = -(input_vector[745] << 7);
assign MEM[5961] = input_vector[745] << 6;
assign MEM[5962] = input_vector[745] << 5;
assign MEM[5963] = input_vector[745] << 4;
assign MEM[5964] = input_vector[745] << 3;
assign MEM[5965] = input_vector[745] << 2;
assign MEM[5966] = input_vector[745] << 1;
assign MEM[5967] = input_vector[745] << 0;
assign MEM[5968] = -(input_vector[746] << 7);
assign MEM[5969] = input_vector[746] << 6;
assign MEM[5970] = input_vector[746] << 5;
assign MEM[5971] = input_vector[746] << 4;
assign MEM[5972] = input_vector[746] << 3;
assign MEM[5973] = input_vector[746] << 2;
assign MEM[5974] = input_vector[746] << 1;
assign MEM[5975] = input_vector[746] << 0;
assign MEM[5976] = -(input_vector[747] << 7);
assign MEM[5977] = input_vector[747] << 6;
assign MEM[5978] = input_vector[747] << 5;
assign MEM[5979] = input_vector[747] << 4;
assign MEM[5980] = input_vector[747] << 3;
assign MEM[5981] = input_vector[747] << 2;
assign MEM[5982] = input_vector[747] << 1;
assign MEM[5983] = input_vector[747] << 0;
assign MEM[5984] = -(input_vector[748] << 7);
assign MEM[5985] = input_vector[748] << 6;
assign MEM[5986] = input_vector[748] << 5;
assign MEM[5987] = input_vector[748] << 4;
assign MEM[5988] = input_vector[748] << 3;
assign MEM[5989] = input_vector[748] << 2;
assign MEM[5990] = input_vector[748] << 1;
assign MEM[5991] = input_vector[748] << 0;
assign MEM[5992] = -(input_vector[749] << 7);
assign MEM[5993] = input_vector[749] << 6;
assign MEM[5994] = input_vector[749] << 5;
assign MEM[5995] = input_vector[749] << 4;
assign MEM[5996] = input_vector[749] << 3;
assign MEM[5997] = input_vector[749] << 2;
assign MEM[5998] = input_vector[749] << 1;
assign MEM[5999] = input_vector[749] << 0;
assign MEM[6000] = -(input_vector[750] << 7);
assign MEM[6001] = input_vector[750] << 6;
assign MEM[6002] = input_vector[750] << 5;
assign MEM[6003] = input_vector[750] << 4;
assign MEM[6004] = input_vector[750] << 3;
assign MEM[6005] = input_vector[750] << 2;
assign MEM[6006] = input_vector[750] << 1;
assign MEM[6007] = input_vector[750] << 0;
assign MEM[6008] = -(input_vector[751] << 7);
assign MEM[6009] = input_vector[751] << 6;
assign MEM[6010] = input_vector[751] << 5;
assign MEM[6011] = input_vector[751] << 4;
assign MEM[6012] = input_vector[751] << 3;
assign MEM[6013] = input_vector[751] << 2;
assign MEM[6014] = input_vector[751] << 1;
assign MEM[6015] = input_vector[751] << 0;
assign MEM[6016] = -(input_vector[752] << 7);
assign MEM[6017] = input_vector[752] << 6;
assign MEM[6018] = input_vector[752] << 5;
assign MEM[6019] = input_vector[752] << 4;
assign MEM[6020] = input_vector[752] << 3;
assign MEM[6021] = input_vector[752] << 2;
assign MEM[6022] = input_vector[752] << 1;
assign MEM[6023] = input_vector[752] << 0;
assign MEM[6024] = -(input_vector[753] << 7);
assign MEM[6025] = input_vector[753] << 6;
assign MEM[6026] = input_vector[753] << 5;
assign MEM[6027] = input_vector[753] << 4;
assign MEM[6028] = input_vector[753] << 3;
assign MEM[6029] = input_vector[753] << 2;
assign MEM[6030] = input_vector[753] << 1;
assign MEM[6031] = input_vector[753] << 0;
assign MEM[6032] = -(input_vector[754] << 7);
assign MEM[6033] = input_vector[754] << 6;
assign MEM[6034] = input_vector[754] << 5;
assign MEM[6035] = input_vector[754] << 4;
assign MEM[6036] = input_vector[754] << 3;
assign MEM[6037] = input_vector[754] << 2;
assign MEM[6038] = input_vector[754] << 1;
assign MEM[6039] = input_vector[754] << 0;
assign MEM[6040] = -(input_vector[755] << 7);
assign MEM[6041] = input_vector[755] << 6;
assign MEM[6042] = input_vector[755] << 5;
assign MEM[6043] = input_vector[755] << 4;
assign MEM[6044] = input_vector[755] << 3;
assign MEM[6045] = input_vector[755] << 2;
assign MEM[6046] = input_vector[755] << 1;
assign MEM[6047] = input_vector[755] << 0;
assign MEM[6048] = -(input_vector[756] << 7);
assign MEM[6049] = input_vector[756] << 6;
assign MEM[6050] = input_vector[756] << 5;
assign MEM[6051] = input_vector[756] << 4;
assign MEM[6052] = input_vector[756] << 3;
assign MEM[6053] = input_vector[756] << 2;
assign MEM[6054] = input_vector[756] << 1;
assign MEM[6055] = input_vector[756] << 0;
assign MEM[6056] = -(input_vector[757] << 7);
assign MEM[6057] = input_vector[757] << 6;
assign MEM[6058] = input_vector[757] << 5;
assign MEM[6059] = input_vector[757] << 4;
assign MEM[6060] = input_vector[757] << 3;
assign MEM[6061] = input_vector[757] << 2;
assign MEM[6062] = input_vector[757] << 1;
assign MEM[6063] = input_vector[757] << 0;
assign MEM[6064] = -(input_vector[758] << 7);
assign MEM[6065] = input_vector[758] << 6;
assign MEM[6066] = input_vector[758] << 5;
assign MEM[6067] = input_vector[758] << 4;
assign MEM[6068] = input_vector[758] << 3;
assign MEM[6069] = input_vector[758] << 2;
assign MEM[6070] = input_vector[758] << 1;
assign MEM[6071] = input_vector[758] << 0;
assign MEM[6072] = -(input_vector[759] << 7);
assign MEM[6073] = input_vector[759] << 6;
assign MEM[6074] = input_vector[759] << 5;
assign MEM[6075] = input_vector[759] << 4;
assign MEM[6076] = input_vector[759] << 3;
assign MEM[6077] = input_vector[759] << 2;
assign MEM[6078] = input_vector[759] << 1;
assign MEM[6079] = input_vector[759] << 0;
assign MEM[6080] = -(input_vector[760] << 7);
assign MEM[6081] = input_vector[760] << 6;
assign MEM[6082] = input_vector[760] << 5;
assign MEM[6083] = input_vector[760] << 4;
assign MEM[6084] = input_vector[760] << 3;
assign MEM[6085] = input_vector[760] << 2;
assign MEM[6086] = input_vector[760] << 1;
assign MEM[6087] = input_vector[760] << 0;
assign MEM[6088] = -(input_vector[761] << 7);
assign MEM[6089] = input_vector[761] << 6;
assign MEM[6090] = input_vector[761] << 5;
assign MEM[6091] = input_vector[761] << 4;
assign MEM[6092] = input_vector[761] << 3;
assign MEM[6093] = input_vector[761] << 2;
assign MEM[6094] = input_vector[761] << 1;
assign MEM[6095] = input_vector[761] << 0;
assign MEM[6096] = -(input_vector[762] << 7);
assign MEM[6097] = input_vector[762] << 6;
assign MEM[6098] = input_vector[762] << 5;
assign MEM[6099] = input_vector[762] << 4;
assign MEM[6100] = input_vector[762] << 3;
assign MEM[6101] = input_vector[762] << 2;
assign MEM[6102] = input_vector[762] << 1;
assign MEM[6103] = input_vector[762] << 0;
assign MEM[6104] = -(input_vector[763] << 7);
assign MEM[6105] = input_vector[763] << 6;
assign MEM[6106] = input_vector[763] << 5;
assign MEM[6107] = input_vector[763] << 4;
assign MEM[6108] = input_vector[763] << 3;
assign MEM[6109] = input_vector[763] << 2;
assign MEM[6110] = input_vector[763] << 1;
assign MEM[6111] = input_vector[763] << 0;
assign MEM[6112] = -(input_vector[764] << 7);
assign MEM[6113] = input_vector[764] << 6;
assign MEM[6114] = input_vector[764] << 5;
assign MEM[6115] = input_vector[764] << 4;
assign MEM[6116] = input_vector[764] << 3;
assign MEM[6117] = input_vector[764] << 2;
assign MEM[6118] = input_vector[764] << 1;
assign MEM[6119] = input_vector[764] << 0;
assign MEM[6120] = -(input_vector[765] << 7);
assign MEM[6121] = input_vector[765] << 6;
assign MEM[6122] = input_vector[765] << 5;
assign MEM[6123] = input_vector[765] << 4;
assign MEM[6124] = input_vector[765] << 3;
assign MEM[6125] = input_vector[765] << 2;
assign MEM[6126] = input_vector[765] << 1;
assign MEM[6127] = input_vector[765] << 0;
assign MEM[6128] = -(input_vector[766] << 7);
assign MEM[6129] = input_vector[766] << 6;
assign MEM[6130] = input_vector[766] << 5;
assign MEM[6131] = input_vector[766] << 4;
assign MEM[6132] = input_vector[766] << 3;
assign MEM[6133] = input_vector[766] << 2;
assign MEM[6134] = input_vector[766] << 1;
assign MEM[6135] = input_vector[766] << 0;
assign MEM[6136] = -(input_vector[767] << 7);
assign MEM[6137] = input_vector[767] << 6;
assign MEM[6138] = input_vector[767] << 5;
assign MEM[6139] = input_vector[767] << 4;
assign MEM[6140] = input_vector[767] << 3;
assign MEM[6141] = input_vector[767] << 2;
assign MEM[6142] = input_vector[767] << 1;
assign MEM[6143] = input_vector[767] << 0;
assign MEM[6144] = -(input_vector[768] << 7);
assign MEM[6145] = input_vector[768] << 6;
assign MEM[6146] = input_vector[768] << 5;
assign MEM[6147] = input_vector[768] << 4;
assign MEM[6148] = input_vector[768] << 3;
assign MEM[6149] = input_vector[768] << 2;
assign MEM[6150] = input_vector[768] << 1;
assign MEM[6151] = input_vector[768] << 0;
assign MEM[6152] = -(input_vector[769] << 7);
assign MEM[6153] = input_vector[769] << 6;
assign MEM[6154] = input_vector[769] << 5;
assign MEM[6155] = input_vector[769] << 4;
assign MEM[6156] = input_vector[769] << 3;
assign MEM[6157] = input_vector[769] << 2;
assign MEM[6158] = input_vector[769] << 1;
assign MEM[6159] = input_vector[769] << 0;
assign MEM[6160] = -(input_vector[770] << 7);
assign MEM[6161] = input_vector[770] << 6;
assign MEM[6162] = input_vector[770] << 5;
assign MEM[6163] = input_vector[770] << 4;
assign MEM[6164] = input_vector[770] << 3;
assign MEM[6165] = input_vector[770] << 2;
assign MEM[6166] = input_vector[770] << 1;
assign MEM[6167] = input_vector[770] << 0;
assign MEM[6168] = -(input_vector[771] << 7);
assign MEM[6169] = input_vector[771] << 6;
assign MEM[6170] = input_vector[771] << 5;
assign MEM[6171] = input_vector[771] << 4;
assign MEM[6172] = input_vector[771] << 3;
assign MEM[6173] = input_vector[771] << 2;
assign MEM[6174] = input_vector[771] << 1;
assign MEM[6175] = input_vector[771] << 0;
assign MEM[6176] = -(input_vector[772] << 7);
assign MEM[6177] = input_vector[772] << 6;
assign MEM[6178] = input_vector[772] << 5;
assign MEM[6179] = input_vector[772] << 4;
assign MEM[6180] = input_vector[772] << 3;
assign MEM[6181] = input_vector[772] << 2;
assign MEM[6182] = input_vector[772] << 1;
assign MEM[6183] = input_vector[772] << 0;
assign MEM[6184] = -(input_vector[773] << 7);
assign MEM[6185] = input_vector[773] << 6;
assign MEM[6186] = input_vector[773] << 5;
assign MEM[6187] = input_vector[773] << 4;
assign MEM[6188] = input_vector[773] << 3;
assign MEM[6189] = input_vector[773] << 2;
assign MEM[6190] = input_vector[773] << 1;
assign MEM[6191] = input_vector[773] << 0;
assign MEM[6192] = -(input_vector[774] << 7);
assign MEM[6193] = input_vector[774] << 6;
assign MEM[6194] = input_vector[774] << 5;
assign MEM[6195] = input_vector[774] << 4;
assign MEM[6196] = input_vector[774] << 3;
assign MEM[6197] = input_vector[774] << 2;
assign MEM[6198] = input_vector[774] << 1;
assign MEM[6199] = input_vector[774] << 0;
assign MEM[6200] = -(input_vector[775] << 7);
assign MEM[6201] = input_vector[775] << 6;
assign MEM[6202] = input_vector[775] << 5;
assign MEM[6203] = input_vector[775] << 4;
assign MEM[6204] = input_vector[775] << 3;
assign MEM[6205] = input_vector[775] << 2;
assign MEM[6206] = input_vector[775] << 1;
assign MEM[6207] = input_vector[775] << 0;
assign MEM[6208] = -(input_vector[776] << 7);
assign MEM[6209] = input_vector[776] << 6;
assign MEM[6210] = input_vector[776] << 5;
assign MEM[6211] = input_vector[776] << 4;
assign MEM[6212] = input_vector[776] << 3;
assign MEM[6213] = input_vector[776] << 2;
assign MEM[6214] = input_vector[776] << 1;
assign MEM[6215] = input_vector[776] << 0;
assign MEM[6216] = -(input_vector[777] << 7);
assign MEM[6217] = input_vector[777] << 6;
assign MEM[6218] = input_vector[777] << 5;
assign MEM[6219] = input_vector[777] << 4;
assign MEM[6220] = input_vector[777] << 3;
assign MEM[6221] = input_vector[777] << 2;
assign MEM[6222] = input_vector[777] << 1;
assign MEM[6223] = input_vector[777] << 0;
assign MEM[6224] = -(input_vector[778] << 7);
assign MEM[6225] = input_vector[778] << 6;
assign MEM[6226] = input_vector[778] << 5;
assign MEM[6227] = input_vector[778] << 4;
assign MEM[6228] = input_vector[778] << 3;
assign MEM[6229] = input_vector[778] << 2;
assign MEM[6230] = input_vector[778] << 1;
assign MEM[6231] = input_vector[778] << 0;
assign MEM[6232] = -(input_vector[779] << 7);
assign MEM[6233] = input_vector[779] << 6;
assign MEM[6234] = input_vector[779] << 5;
assign MEM[6235] = input_vector[779] << 4;
assign MEM[6236] = input_vector[779] << 3;
assign MEM[6237] = input_vector[779] << 2;
assign MEM[6238] = input_vector[779] << 1;
assign MEM[6239] = input_vector[779] << 0;
assign MEM[6240] = -(input_vector[780] << 7);
assign MEM[6241] = input_vector[780] << 6;
assign MEM[6242] = input_vector[780] << 5;
assign MEM[6243] = input_vector[780] << 4;
assign MEM[6244] = input_vector[780] << 3;
assign MEM[6245] = input_vector[780] << 2;
assign MEM[6246] = input_vector[780] << 1;
assign MEM[6247] = input_vector[780] << 0;
assign MEM[6248] = -(input_vector[781] << 7);
assign MEM[6249] = input_vector[781] << 6;
assign MEM[6250] = input_vector[781] << 5;
assign MEM[6251] = input_vector[781] << 4;
assign MEM[6252] = input_vector[781] << 3;
assign MEM[6253] = input_vector[781] << 2;
assign MEM[6254] = input_vector[781] << 1;
assign MEM[6255] = input_vector[781] << 0;
assign MEM[6256] = -(input_vector[782] << 7);
assign MEM[6257] = input_vector[782] << 6;
assign MEM[6258] = input_vector[782] << 5;
assign MEM[6259] = input_vector[782] << 4;
assign MEM[6260] = input_vector[782] << 3;
assign MEM[6261] = input_vector[782] << 2;
assign MEM[6262] = input_vector[782] << 1;
assign MEM[6263] = input_vector[782] << 0;
assign MEM[6264] = -(input_vector[783] << 7);
assign MEM[6265] = input_vector[783] << 6;
assign MEM[6266] = input_vector[783] << 5;
assign MEM[6267] = input_vector[783] << 4;
assign MEM[6268] = input_vector[783] << 3;
assign MEM[6269] = input_vector[783] << 2;
assign MEM[6270] = input_vector[783] << 1;
assign MEM[6271] = input_vector[783] << 0;
assign MEM[6272] = MEM[3384] + MEM[3385];
assign MEM[6273] = MEM[4752] + MEM[4753];
assign MEM[6274] = MEM[1072] + MEM[1073];
assign MEM[6275] = MEM[2280] + MEM[2281];
assign MEM[6276] = MEM[3616] + MEM[3617];
assign MEM[6277] = MEM[4113] + MEM[4112];
assign MEM[6278] = MEM[6120] + MEM[6121];
assign MEM[6279] = MEM[6122] + MEM[6278];
assign MEM[6280] = MEM[304] + MEM[305];
assign MEM[6281] = MEM[1064] + MEM[1065];
assign MEM[6282] = MEM[2496] + MEM[2497];
assign MEM[6283] = MEM[2816] + MEM[2817];
assign MEM[6284] = MEM[3624] + MEM[3625];
assign MEM[6285] = MEM[3744] + MEM[3745];
assign MEM[6286] = MEM[4448] + MEM[4449];
assign MEM[6287] = MEM[6280] + MEM[306];
assign MEM[6288] = MEM[1761] + MEM[1760];
assign MEM[6289] = MEM[2729] + MEM[2728];
assign MEM[6290] = MEM[2936] + MEM[2937];
assign MEM[6291] = MEM[2953] + MEM[2952];
assign MEM[6292] = MEM[3128] + MEM[3129];
assign MEM[6293] = MEM[3288] + MEM[3289];
assign MEM[6294] = MEM[3736] + MEM[3737];
assign MEM[6295] = MEM[3984] + MEM[3985];
assign MEM[6296] = MEM[4072] + MEM[4073];
assign MEM[6297] = MEM[4105] + MEM[4104];
assign MEM[6298] = MEM[4304] + MEM[4305];
assign MEM[6299] = MEM[4344] + MEM[4345];
assign MEM[6300] = MEM[4744] + MEM[4745];
assign MEM[6301] = MEM[5193] + MEM[5192];
assign MEM[6302] = MEM[6292] + MEM[3130];
assign MEM[6303] = MEM[528] + MEM[529];
assign MEM[6304] = MEM[1288] + MEM[1289];
assign MEM[6305] = MEM[1832] + MEM[1833];
assign MEM[6306] = MEM[2480] + MEM[2481];
assign MEM[6307] = MEM[3312] + MEM[3313];
assign MEM[6308] = MEM[3728] + MEM[3729];
assign MEM[6309] = MEM[3848] + MEM[3849];
assign MEM[6310] = MEM[3968] + MEM[3969];
assign MEM[6311] = MEM[3977] + MEM[3976];
assign MEM[6312] = MEM[4088] + MEM[4089];
assign MEM[6313] = MEM[4097] + MEM[4096];
assign MEM[6314] = MEM[4152] + MEM[4153];
assign MEM[6315] = MEM[4296] + MEM[4297];
assign MEM[6316] = MEM[5360] + MEM[5361];
assign MEM[6317] = MEM[5362] + MEM[6316];
assign MEM[6318] = MEM[5776] + MEM[5777];
assign MEM[6319] = MEM[232] + MEM[233];
assign MEM[6320] = MEM[234] + MEM[235];
assign MEM[6321] = MEM[236] + MEM[6319];
assign MEM[6322] = MEM[328] + MEM[329];
assign MEM[6323] = MEM[552] + MEM[553];
assign MEM[6324] = MEM[1056] + MEM[1057];
assign MEM[6325] = MEM[1160] + MEM[1161];
assign MEM[6326] = MEM[2056] + MEM[2057];
assign MEM[6327] = MEM[2361] + MEM[2360];
assign MEM[6328] = MEM[2504] + MEM[2505];
assign MEM[6329] = MEM[2545] + MEM[2544];
assign MEM[6330] = MEM[2561] + MEM[2560];
assign MEM[6331] = MEM[2585] + MEM[2584];
assign MEM[6332] = MEM[2753] + MEM[2752];
assign MEM[6333] = MEM[2840] + MEM[2841];
assign MEM[6334] = MEM[2888] + MEM[2889];
assign MEM[6335] = MEM[3064] + MEM[3065];
assign MEM[6336] = MEM[3089] + MEM[3088];
assign MEM[6337] = MEM[3112] + MEM[3113];
assign MEM[6338] = MEM[3336] + MEM[3337];
assign MEM[6339] = MEM[3512] + MEM[3513];
assign MEM[6340] = MEM[3520] + MEM[3521];
assign MEM[6341] = MEM[3840] + MEM[3841];
assign MEM[6342] = MEM[3881] + MEM[3880];
assign MEM[6343] = MEM[4216] + MEM[4217];
assign MEM[6344] = MEM[4336] + MEM[4337];
assign MEM[6345] = MEM[4648] + MEM[4649];
assign MEM[6346] = MEM[5416] + MEM[5417];
assign MEM[6347] = MEM[5552] + MEM[5553];
assign MEM[6348] = MEM[6320] + MEM[6321];
assign MEM[6349] = MEM[200] + MEM[201];
assign MEM[6350] = MEM[202] + MEM[203];
assign MEM[6351] = MEM[204] + MEM[6349];
assign MEM[6352] = MEM[288] + MEM[289];
assign MEM[6353] = MEM[290] + MEM[6352];
assign MEM[6354] = MEM[352] + MEM[353];
assign MEM[6355] = MEM[440] + MEM[441];
assign MEM[6356] = MEM[442] + MEM[443];
assign MEM[6357] = MEM[444] + MEM[6355];
assign MEM[6358] = MEM[512] + MEM[513];
assign MEM[6359] = MEM[808] + MEM[809];
assign MEM[6360] = MEM[1080] + MEM[1081];
assign MEM[6361] = MEM[1297] + MEM[1296];
assign MEM[6362] = MEM[1616] + MEM[1617];
assign MEM[6363] = MEM[2345] + MEM[2344];
assign MEM[6364] = MEM[2568] + MEM[2569];
assign MEM[6365] = MEM[2576] + MEM[2577];
assign MEM[6366] = MEM[2641] + MEM[2640];
assign MEM[6367] = MEM[2744] + MEM[2745];
assign MEM[6368] = MEM[2769] + MEM[2768];
assign MEM[6369] = MEM[2857] + MEM[2856];
assign MEM[6370] = MEM[2865] + MEM[2864];
assign MEM[6371] = MEM[2896] + MEM[2897];
assign MEM[6372] = MEM[2945] + MEM[2944];
assign MEM[6373] = MEM[2976] + MEM[2977];
assign MEM[6374] = MEM[3072] + MEM[3073];
assign MEM[6375] = MEM[3321] + MEM[3320];
assign MEM[6376] = MEM[3328] + MEM[3329];
assign MEM[6377] = MEM[3496] + MEM[3497];
assign MEM[6378] = MEM[3992] + MEM[3993];
assign MEM[6379] = MEM[4121] + MEM[4120];
assign MEM[6380] = MEM[4496] + MEM[4497];
assign MEM[6381] = MEM[4672] + MEM[4673];
assign MEM[6382] = MEM[4920] + MEM[4921];
assign MEM[6383] = MEM[4922] + MEM[4923];
assign MEM[6384] = MEM[4924] + MEM[6382];
assign MEM[6385] = MEM[5320] + MEM[5321];
assign MEM[6386] = MEM[5528] + MEM[5529];
assign MEM[6387] = MEM[6224] + MEM[6225];
assign MEM[6388] = MEM[6226] + MEM[6387];
assign MEM[6389] = MEM[6350] + MEM[6351];
assign MEM[6390] = MEM[6356] + MEM[6357];
assign MEM[6391] = MEM[6383] + MEM[6384];
assign MEM[6392] = MEM[96] + MEM[97];
assign MEM[6393] = MEM[98] + MEM[99];
assign MEM[6394] = MEM[100] + MEM[6392];
assign MEM[6395] = MEM[224] + MEM[225];
assign MEM[6396] = MEM[226] + MEM[227];
assign MEM[6397] = MEM[228] + MEM[6395];
assign MEM[6398] = MEM[248] + MEM[249];
assign MEM[6399] = MEM[250] + MEM[251];
assign MEM[6400] = MEM[252] + MEM[6398];
assign MEM[6401] = MEM[296] + MEM[297];
assign MEM[6402] = MEM[298] + MEM[6401];
assign MEM[6403] = MEM[912] + MEM[913];
assign MEM[6404] = MEM[914] + MEM[6403];
assign MEM[6405] = MEM[936] + MEM[937];
assign MEM[6406] = MEM[1128] + MEM[1129];
assign MEM[6407] = MEM[1130] + MEM[1131];
assign MEM[6408] = MEM[1132] + MEM[6406];
assign MEM[6409] = MEM[1240] + MEM[1241];
assign MEM[6410] = MEM[1400] + MEM[1401];
assign MEM[6411] = MEM[1424] + MEM[1425];
assign MEM[6412] = MEM[1488] + MEM[1489];
assign MEM[6413] = MEM[1496] + MEM[1497];
assign MEM[6414] = MEM[1504] + MEM[1505];
assign MEM[6415] = MEM[1512] + MEM[1513];
assign MEM[6416] = MEM[1624] + MEM[1625];
assign MEM[6417] = MEM[1840] + MEM[1841];
assign MEM[6418] = MEM[1977] + MEM[1976];
assign MEM[6419] = MEM[2032] + MEM[2033];
assign MEM[6420] = MEM[2104] + MEM[2105];
assign MEM[6421] = MEM[2537] + MEM[2536];
assign MEM[6422] = MEM[2649] + MEM[2648];
assign MEM[6423] = MEM[3096] + MEM[3097];
assign MEM[6424] = MEM[3208] + MEM[3209];
assign MEM[6425] = MEM[3865] + MEM[3864];
assign MEM[6426] = MEM[3888] + MEM[3889];
assign MEM[6427] = MEM[3952] + MEM[3953];
assign MEM[6428] = MEM[3960] + MEM[3961];
assign MEM[6429] = MEM[4064] + MEM[4065];
assign MEM[6430] = MEM[4154] + MEM[6314];
assign MEM[6431] = MEM[4632] + MEM[4633];
assign MEM[6432] = MEM[4832] + MEM[4833];
assign MEM[6433] = MEM[4864] + MEM[4865];
assign MEM[6434] = MEM[4872] + MEM[4873];
assign MEM[6435] = MEM[5072] + MEM[5073];
assign MEM[6436] = MEM[5120] + MEM[5121];
assign MEM[6437] = MEM[5168] + MEM[5169];
assign MEM[6438] = MEM[5170] + MEM[6437];
assign MEM[6439] = MEM[5200] + MEM[5201];
assign MEM[6440] = MEM[5352] + MEM[5353];
assign MEM[6441] = MEM[5632] + MEM[5633];
assign MEM[6442] = MEM[6152] + MEM[6153];
assign MEM[6443] = MEM[6393] + MEM[6394];
assign MEM[6444] = MEM[6396] + MEM[6397];
assign MEM[6445] = MEM[6399] + MEM[6400];
assign MEM[6446] = MEM[6407] + MEM[6408];
assign MEM[6447] = MEM[216] + MEM[217];
assign MEM[6448] = MEM[218] + MEM[219];
assign MEM[6449] = MEM[220] + MEM[6447];
assign MEM[6450] = MEM[264] + MEM[265];
assign MEM[6451] = MEM[266] + MEM[267];
assign MEM[6452] = MEM[268] + MEM[6450];
assign MEM[6453] = MEM[536] + MEM[537];
assign MEM[6454] = MEM[648] + MEM[649];
assign MEM[6455] = MEM[650] + MEM[6454];
assign MEM[6456] = MEM[672] + MEM[673];
assign MEM[6457] = MEM[674] + MEM[675];
assign MEM[6458] = MEM[676] + MEM[6456];
assign MEM[6459] = MEM[680] + MEM[681];
assign MEM[6460] = MEM[682] + MEM[683];
assign MEM[6461] = MEM[684] + MEM[6459];
assign MEM[6462] = MEM[729] + MEM[728];
assign MEM[6463] = MEM[768] + MEM[769];
assign MEM[6464] = MEM[792] + MEM[793];
assign MEM[6465] = MEM[872] + MEM[873];
assign MEM[6466] = MEM[1416] + MEM[1417];
assign MEM[6467] = MEM[1440] + MEM[1441];
assign MEM[6468] = MEM[1521] + MEM[1520];
assign MEM[6469] = MEM[1784] + MEM[1785];
assign MEM[6470] = MEM[1786] + MEM[6469];
assign MEM[6471] = MEM[1872] + MEM[1873];
assign MEM[6472] = MEM[1952] + MEM[1953];
assign MEM[6473] = MEM[2417] + MEM[2416];
assign MEM[6474] = MEM[2425] + MEM[2424];
assign MEM[6475] = MEM[2472] + MEM[2473];
assign MEM[6476] = MEM[2474] + MEM[6475];
assign MEM[6477] = MEM[2488] + MEM[2489];
assign MEM[6478] = MEM[2633] + MEM[2632];
assign MEM[6479] = MEM[2696] + MEM[2697];
assign MEM[6480] = MEM[2698] + MEM[6479];
assign MEM[6481] = MEM[2881] + MEM[2880];
assign MEM[6482] = MEM[2920] + MEM[2921];
assign MEM[6483] = MEM[2922] + MEM[2923];
assign MEM[6484] = MEM[2985] + MEM[2984];
assign MEM[6485] = MEM[3120] + MEM[3121];
assign MEM[6486] = MEM[3169] + MEM[3168];
assign MEM[6487] = MEM[3344] + MEM[3345];
assign MEM[6488] = MEM[3400] + MEM[3401];
assign MEM[6489] = MEM[3488] + MEM[3489];
assign MEM[6490] = MEM[3499] + MEM[503];
assign MEM[6491] = MEM[3576] + MEM[3577];
assign MEM[6492] = MEM[3657] + MEM[3656];
assign MEM[6493] = MEM[3752] + MEM[3753];
assign MEM[6494] = MEM[3944] + MEM[3945];
assign MEM[6495] = MEM[4080] + MEM[4081];
assign MEM[6496] = MEM[4129] + MEM[4128];
assign MEM[6497] = MEM[4200] + MEM[4201];
assign MEM[6498] = MEM[4320] + MEM[4321];
assign MEM[6499] = MEM[4529] + MEM[4528];
assign MEM[6500] = MEM[4834] + MEM[6432];
assign MEM[6501] = MEM[5297] + MEM[5296];
assign MEM[6502] = MEM[5816] + MEM[5817];
assign MEM[6503] = MEM[5818] + MEM[5819];
assign MEM[6504] = MEM[5820] + MEM[6502];
assign MEM[6505] = MEM[5872] + MEM[5873];
assign MEM[6506] = MEM[5913] + MEM[5912];
assign MEM[6507] = MEM[6000] + MEM[6001];
assign MEM[6508] = MEM[6016] + MEM[6017];
assign MEM[6509] = MEM[6018] + MEM[6019];
assign MEM[6510] = MEM[6020] + MEM[6508];
assign MEM[6511] = MEM[6200] + MEM[6201];
assign MEM[6512] = MEM[6202] + MEM[6511];
assign MEM[6513] = MEM[6448] + MEM[6449];
assign MEM[6514] = MEM[6451] + MEM[6452];
assign MEM[6515] = MEM[6457] + MEM[6458];
assign MEM[6516] = MEM[6460] + MEM[6461];
assign MEM[6517] = MEM[6482] + MEM[6483];
assign MEM[6518] = MEM[6503] + MEM[6504];
assign MEM[6519] = MEM[6509] + MEM[6510];
assign MEM[6520] = MEM[72] + MEM[73];
assign MEM[6521] = MEM[74] + MEM[75];
assign MEM[6522] = MEM[76] + MEM[6520];
assign MEM[6523] = MEM[149] + MEM[990];
assign MEM[6524] = MEM[336] + MEM[337];
assign MEM[6525] = MEM[397] + MEM[1211];
assign MEM[6526] = MEM[424] + MEM[425];
assign MEM[6527] = MEM[426] + MEM[427];
assign MEM[6528] = MEM[428] + MEM[6526];
assign MEM[6529] = MEM[432] + MEM[433];
assign MEM[6530] = MEM[434] + MEM[435];
assign MEM[6531] = MEM[436] + MEM[6529];
assign MEM[6532] = MEM[462] + MEM[2363];
assign MEM[6533] = MEM[496] + MEM[497];
assign MEM[6534] = MEM[498] + MEM[6533];
assign MEM[6535] = MEM[504] + MEM[505];
assign MEM[6536] = MEM[544] + MEM[545];
assign MEM[6537] = MEM[824] + MEM[825];
assign MEM[6538] = MEM[848] + MEM[849];
assign MEM[6539] = MEM[888] + MEM[889];
assign MEM[6540] = MEM[890] + MEM[891];
assign MEM[6541] = MEM[892] + MEM[6539];
assign MEM[6542] = MEM[920] + MEM[921];
assign MEM[6543] = MEM[922] + MEM[923];
assign MEM[6544] = MEM[924] + MEM[6542];
assign MEM[6545] = MEM[1088] + MEM[1089];
assign MEM[6546] = MEM[1168] + MEM[1169];
assign MEM[6547] = MEM[1208] + MEM[1209];
assign MEM[6548] = MEM[1280] + MEM[1281];
assign MEM[6549] = MEM[1336] + MEM[1337];
assign MEM[6550] = MEM[1338] + MEM[1339];
assign MEM[6551] = MEM[1340] + MEM[6549];
assign MEM[6552] = MEM[1352] + MEM[1353];
assign MEM[6553] = MEM[1354] + MEM[1355];
assign MEM[6554] = MEM[1356] + MEM[6552];
assign MEM[6555] = MEM[1574] + MEM[2791];
assign MEM[6556] = MEM[1729] + MEM[1728];
assign MEM[6557] = MEM[1808] + MEM[1809];
assign MEM[6558] = MEM[1842] + MEM[6417];
assign MEM[6559] = MEM[1864] + MEM[1865];
assign MEM[6560] = MEM[2120] + MEM[2121];
assign MEM[6561] = MEM[2192] + MEM[2193];
assign MEM[6562] = MEM[2256] + MEM[2257];
assign MEM[6563] = MEM[2337] + MEM[2336];
assign MEM[6564] = MEM[2512] + MEM[2513];
assign MEM[6565] = MEM[2529] + MEM[2528];
assign MEM[6566] = MEM[2721] + MEM[2720];
assign MEM[6567] = MEM[2737] + MEM[2736];
assign MEM[6568] = MEM[2761] + MEM[2760];
assign MEM[6569] = MEM[2801] + MEM[2800];
assign MEM[6570] = MEM[2961] + MEM[2960];
assign MEM[6571] = MEM[3056] + MEM[3057];
assign MEM[6572] = MEM[3144] + MEM[3145];
assign MEM[6573] = MEM[3146] + MEM[3147];
assign MEM[6574] = MEM[3148] + MEM[6572];
assign MEM[6575] = MEM[3272] + MEM[3273];
assign MEM[6576] = MEM[3392] + MEM[3393];
assign MEM[6577] = MEM[3448] + MEM[3449];
assign MEM[6578] = MEM[3528] + MEM[3529];
assign MEM[6579] = MEM[3560] + MEM[3561];
assign MEM[6580] = MEM[3633] + MEM[3632];
assign MEM[6581] = MEM[3641] + MEM[3640];
assign MEM[6582] = MEM[3649] + MEM[3648];
assign MEM[6583] = MEM[3680] + MEM[3681];
assign MEM[6584] = MEM[3704] + MEM[3705];
assign MEM[6585] = MEM[3857] + MEM[3856];
assign MEM[6586] = MEM[3873] + MEM[3872];
assign MEM[6587] = MEM[4168] + MEM[4169];
assign MEM[6588] = MEM[4312] + MEM[4313];
assign MEM[6589] = MEM[4641] + MEM[4640];
assign MEM[6590] = MEM[4664] + MEM[4665];
assign MEM[6591] = MEM[4969] + MEM[4968];
assign MEM[6592] = MEM[5112] + MEM[5113];
assign MEM[6593] = MEM[5305] + MEM[5304];
assign MEM[6594] = MEM[5600] + MEM[5601];
assign MEM[6595] = MEM[5602] + MEM[5603];
assign MEM[6596] = MEM[5604] + MEM[6594];
assign MEM[6597] = MEM[5640] + MEM[5641];
assign MEM[6598] = MEM[5760] + MEM[5761];
assign MEM[6599] = MEM[5800] + MEM[5801];
assign MEM[6600] = MEM[5802] + MEM[5803];
assign MEM[6601] = MEM[5804] + MEM[6599];
assign MEM[6602] = MEM[5840] + MEM[5841];
assign MEM[6603] = MEM[5842] + MEM[5843];
assign MEM[6604] = MEM[5844] + MEM[6602];
assign MEM[6605] = MEM[5960] + MEM[5961];
assign MEM[6606] = MEM[6168] + MEM[6169];
assign MEM[6607] = MEM[6216] + MEM[6217];
assign MEM[6608] = MEM[6218] + MEM[6607];
assign MEM[6609] = MEM[6521] + MEM[6522];
assign MEM[6610] = MEM[6527] + MEM[6528];
assign MEM[6611] = MEM[6530] + MEM[6531];
assign MEM[6612] = MEM[6535] + MEM[506];
assign MEM[6613] = MEM[6540] + MEM[6541];
assign MEM[6614] = MEM[6543] + MEM[6544];
assign MEM[6615] = MEM[6550] + MEM[6551];
assign MEM[6616] = MEM[6553] + MEM[6554];
assign MEM[6617] = MEM[6573] + MEM[6574];
assign MEM[6618] = MEM[6595] + MEM[6596];
assign MEM[6619] = MEM[6600] + MEM[6601];
assign MEM[6620] = MEM[6603] + MEM[6604];
assign MEM[6621] = MEM[160] + MEM[161];
assign MEM[6622] = MEM[162] + MEM[163];
assign MEM[6623] = MEM[164] + MEM[6621];
assign MEM[6624] = MEM[192] + MEM[193];
assign MEM[6625] = MEM[194] + MEM[195];
assign MEM[6626] = MEM[196] + MEM[6624];
assign MEM[6627] = MEM[272] + MEM[273];
assign MEM[6628] = MEM[274] + MEM[275];
assign MEM[6629] = MEM[308] + MEM[2149];
assign MEM[6630] = MEM[344] + MEM[345];
assign MEM[6631] = MEM[368] + MEM[369];
assign MEM[6632] = MEM[384] + MEM[385];
assign MEM[6633] = MEM[540] + MEM[695];
assign MEM[6634] = MEM[568] + MEM[569];
assign MEM[6635] = MEM[724] + MEM[3558];
assign MEM[6636] = MEM[736] + MEM[737];
assign MEM[6637] = MEM[856] + MEM[857];
assign MEM[6638] = MEM[880] + MEM[881];
assign MEM[6639] = MEM[882] + MEM[883];
assign MEM[6640] = MEM[884] + MEM[6638];
assign MEM[6641] = MEM[896] + MEM[897];
assign MEM[6642] = MEM[898] + MEM[899];
assign MEM[6643] = MEM[900] + MEM[6641];
assign MEM[6644] = MEM[944] + MEM[945];
assign MEM[6645] = MEM[1136] + MEM[1137];
assign MEM[6646] = MEM[1138] + MEM[1139];
assign MEM[6647] = MEM[1140] + MEM[6645];
assign MEM[6648] = MEM[1392] + MEM[1393];
assign MEM[6649] = MEM[1418] + MEM[6466];
assign MEM[6650] = MEM[1456] + MEM[1457];
assign MEM[6651] = MEM[1464] + MEM[1465];
assign MEM[6652] = MEM[1524] + MEM[2651];
assign MEM[6653] = MEM[1568] + MEM[1569];
assign MEM[6654] = MEM[1570] + MEM[1571];
assign MEM[6655] = MEM[1572] + MEM[6653];
assign MEM[6656] = MEM[1592] + MEM[1593];
assign MEM[6657] = MEM[1753] + MEM[1752];
assign MEM[6658] = MEM[1866] + MEM[6559];
assign MEM[6659] = MEM[1900] + MEM[4450];
assign MEM[6660] = MEM[1969] + MEM[1968];
assign MEM[6661] = MEM[2110] + MEM[3346];
assign MEM[6662] = MEM[2112] + MEM[2113];
assign MEM[6663] = MEM[2129] + MEM[2128];
assign MEM[6664] = MEM[2232] + MEM[2233];
assign MEM[6665] = MEM[2248] + MEM[2249];
assign MEM[6666] = MEM[2250] + MEM[2251];
assign MEM[6667] = MEM[2353] + MEM[2352];
assign MEM[6668] = MEM[2368] + MEM[2369];
assign MEM[6669] = MEM[2440] + MEM[2441];
assign MEM[6670] = MEM[2461] + MEM[375];
assign MEM[6671] = MEM[2592] + MEM[2593];
assign MEM[6672] = MEM[2704] + MEM[2705];
assign MEM[6673] = MEM[2809] + MEM[2808];
assign MEM[6674] = MEM[2843] + MEM[2943];
assign MEM[6675] = MEM[2873] + MEM[2872];
assign MEM[6676] = MEM[3000] + MEM[3001];
assign MEM[6677] = MEM[3193] + MEM[3192];
assign MEM[6678] = MEM[3224] + MEM[3225];
assign MEM[6679] = MEM[3280] + MEM[3281];
assign MEM[6680] = MEM[3368] + MEM[3369];
assign MEM[6681] = MEM[3391] + MEM[2596];
assign MEM[6682] = MEM[3462] + MEM[2938];
assign MEM[6683] = MEM[3472] + MEM[3473];
assign MEM[6684] = MEM[3504] + MEM[3505];
assign MEM[6685] = MEM[3536] + MEM[3537];
assign MEM[6686] = MEM[3552] + MEM[3553];
assign MEM[6687] = MEM[3584] + MEM[3585];
assign MEM[6688] = MEM[3586] + MEM[3587];
assign MEM[6689] = MEM[3588] + MEM[6687];
assign MEM[6690] = MEM[3608] + MEM[3609];
assign MEM[6691] = MEM[3659] + MEM[1069];
assign MEM[6692] = MEM[3741] + MEM[3311];
assign MEM[6693] = MEM[3792] + MEM[3793];
assign MEM[6694] = MEM[3891] + MEM[396];
assign MEM[6695] = MEM[3905] + MEM[3904];
assign MEM[6696] = MEM[3920] + MEM[3921];
assign MEM[6697] = MEM[3928] + MEM[3929];
assign MEM[6698] = MEM[4000] + MEM[4001];
assign MEM[6699] = MEM[4328] + MEM[4329];
assign MEM[6700] = MEM[4384] + MEM[4385];
assign MEM[6701] = MEM[4416] + MEM[4417];
assign MEM[6702] = MEM[4432] + MEM[4433];
assign MEM[6703] = MEM[4439] + MEM[533];
assign MEM[6704] = MEM[4552] + MEM[4553];
assign MEM[6705] = MEM[4656] + MEM[4657];
assign MEM[6706] = MEM[4760] + MEM[4761];
assign MEM[6707] = MEM[4808] + MEM[4809];
assign MEM[6708] = MEM[4816] + MEM[4817];
assign MEM[6709] = MEM[4848] + MEM[4849];
assign MEM[6710] = MEM[4977] + MEM[4976];
assign MEM[6711] = MEM[5144] + MEM[5145];
assign MEM[6712] = MEM[5146] + MEM[5147];
assign MEM[6713] = MEM[5148] + MEM[6711];
assign MEM[6714] = MEM[5288] + MEM[5289];
assign MEM[6715] = MEM[5613] + MEM[5287];
assign MEM[6716] = MEM[5768] + MEM[5769];
assign MEM[6717] = MEM[5784] + MEM[5785];
assign MEM[6718] = MEM[5815] + MEM[1287];
assign MEM[6719] = MEM[5832] + MEM[5833];
assign MEM[6720] = MEM[5834] + MEM[5835];
assign MEM[6721] = MEM[5836] + MEM[6719];
assign MEM[6722] = MEM[5856] + MEM[5857];
assign MEM[6723] = MEM[5880] + MEM[5881];
assign MEM[6724] = MEM[5888] + MEM[5889];
assign MEM[6725] = MEM[5945] + MEM[5944];
assign MEM[6726] = MEM[6088] + MEM[6089];
assign MEM[6727] = MEM[6090] + MEM[6091];
assign MEM[6728] = MEM[6092] + MEM[6726];
assign MEM[6729] = MEM[6128] + MEM[6129];
assign MEM[6730] = MEM[6232] + MEM[6233];
assign MEM[6731] = MEM[6234] + MEM[6235];
assign MEM[6732] = MEM[6236] + MEM[6730];
assign MEM[6733] = MEM[6248] + MEM[6249];
assign MEM[6734] = MEM[6250] + MEM[6251];
assign MEM[6735] = MEM[6252] + MEM[6733];
assign MEM[6736] = MEM[6276] + MEM[6284];
assign MEM[6737] = MEM[6305] + MEM[1834];
assign MEM[6738] = MEM[6622] + MEM[6623];
assign MEM[6739] = MEM[6625] + MEM[6626];
assign MEM[6740] = MEM[6627] + MEM[6628];
assign MEM[6741] = MEM[6630] + MEM[346];
assign MEM[6742] = MEM[6632] + MEM[386];
assign MEM[6743] = MEM[6639] + MEM[6640];
assign MEM[6744] = MEM[6642] + MEM[6643];
assign MEM[6745] = MEM[6646] + MEM[6647];
assign MEM[6746] = MEM[6654] + MEM[6655];
assign MEM[6747] = MEM[6665] + MEM[6666];
assign MEM[6748] = MEM[6680] + MEM[3370];
assign MEM[6749] = MEM[6688] + MEM[6689];
assign MEM[6750] = MEM[6690] + MEM[3610];
assign MEM[6751] = MEM[6712] + MEM[6713];
assign MEM[6752] = MEM[6720] + MEM[6721];
assign MEM[6753] = MEM[6727] + MEM[6728];
assign MEM[6754] = MEM[6731] + MEM[6732];
assign MEM[6755] = MEM[6734] + MEM[6735];
assign MEM[6756] = MEM[8] + MEM[9];
assign MEM[6757] = MEM[10] + MEM[11];
assign MEM[6758] = MEM[12] + MEM[6756];
assign MEM[6759] = MEM[88] + MEM[89];
assign MEM[6760] = MEM[90] + MEM[91];
assign MEM[6761] = MEM[92] + MEM[6759];
assign MEM[6762] = MEM[120] + MEM[121];
assign MEM[6763] = MEM[122] + MEM[123];
assign MEM[6764] = MEM[124] + MEM[6762];
assign MEM[6765] = MEM[144] + MEM[145];
assign MEM[6766] = MEM[146] + MEM[147];
assign MEM[6767] = MEM[148] + MEM[6765];
assign MEM[6768] = MEM[152] + MEM[153];
assign MEM[6769] = MEM[154] + MEM[155];
assign MEM[6770] = MEM[156] + MEM[6768];
assign MEM[6771] = MEM[168] + MEM[169];
assign MEM[6772] = MEM[170] + MEM[171];
assign MEM[6773] = MEM[172] + MEM[6771];
assign MEM[6774] = MEM[269] + MEM[1006];
assign MEM[6775] = MEM[330] + MEM[1094];
assign MEM[6776] = MEM[360] + MEM[361];
assign MEM[6777] = MEM[392] + MEM[393];
assign MEM[6778] = MEM[394] + MEM[6777];
assign MEM[6779] = MEM[398] + MEM[652];
assign MEM[6780] = MEM[456] + MEM[457];
assign MEM[6781] = MEM[458] + MEM[459];
assign MEM[6782] = MEM[460] + MEM[6780];
assign MEM[6783] = MEM[480] + MEM[481];
assign MEM[6784] = MEM[576] + MEM[577];
assign MEM[6785] = MEM[606] + MEM[2823];
assign MEM[6786] = MEM[640] + MEM[641];
assign MEM[6787] = MEM[642] + MEM[6786];
assign MEM[6788] = MEM[656] + MEM[657];
assign MEM[6789] = MEM[658] + MEM[659];
assign MEM[6790] = MEM[660] + MEM[6788];
assign MEM[6791] = MEM[696] + MEM[697];
assign MEM[6792] = MEM[698] + MEM[699];
assign MEM[6793] = MEM[700] + MEM[6791];
assign MEM[6794] = MEM[712] + MEM[713];
assign MEM[6795] = MEM[714] + MEM[6794];
assign MEM[6796] = MEM[841] + MEM[840];
assign MEM[6797] = MEM[953] + MEM[952];
assign MEM[6798] = MEM[961] + MEM[960];
assign MEM[6799] = MEM[1032] + MEM[1033];
assign MEM[6800] = MEM[1192] + MEM[1193];
assign MEM[6801] = MEM[1197] + MEM[3950];
assign MEM[6802] = MEM[1384] + MEM[1385];
assign MEM[6803] = MEM[1408] + MEM[1409];
assign MEM[6804] = MEM[1608] + MEM[1609];
assign MEM[6805] = MEM[1645] + MEM[2282];
assign MEM[6806] = MEM[1648] + MEM[1649];
assign MEM[6807] = MEM[1672] + MEM[1673];
assign MEM[6808] = MEM[1725] + MEM[1327];
assign MEM[6809] = MEM[1768] + MEM[1769];
assign MEM[6810] = MEM[1771] + MEM[703];
assign MEM[6811] = MEM[1800] + MEM[1801];
assign MEM[6812] = MEM[1802] + MEM[6811];
assign MEM[6813] = MEM[2015] + MEM[4754];
assign MEM[6814] = MEM[2040] + MEM[2041];
assign MEM[6815] = MEM[2132] + MEM[2666];
assign MEM[6816] = MEM[2137] + MEM[2136];
assign MEM[6817] = MEM[2184] + MEM[2185];
assign MEM[6818] = MEM[2321] + MEM[2320];
assign MEM[6819] = MEM[2393] + MEM[2392];
assign MEM[6820] = MEM[2409] + MEM[2408];
assign MEM[6821] = MEM[2552] + MEM[2553];
assign MEM[6822] = MEM[2712] + MEM[2713];
assign MEM[6823] = MEM[2785] + MEM[2784];
assign MEM[6824] = MEM[2904] + MEM[2905];
assign MEM[6825] = MEM[2906] + MEM[2907];
assign MEM[6826] = MEM[2928] + MEM[2929];
assign MEM[6827] = MEM[2969] + MEM[2968];
assign MEM[6828] = MEM[3009] + MEM[3008];
assign MEM[6829] = MEM[3048] + MEM[3049];
assign MEM[6830] = MEM[3075] + MEM[3074];
assign MEM[6831] = MEM[3080] + MEM[3081];
assign MEM[6832] = MEM[3105] + MEM[3104];
assign MEM[6833] = MEM[3136] + MEM[3137];
assign MEM[6834] = MEM[3138] + MEM[3139];
assign MEM[6835] = MEM[3140] + MEM[6833];
assign MEM[6836] = MEM[3160] + MEM[3161];
assign MEM[6837] = MEM[3282] + MEM[6679];
assign MEM[6838] = MEM[3296] + MEM[3297];
assign MEM[6839] = MEM[3409] + MEM[3408];
assign MEM[6840] = MEM[3417] + MEM[3416];
assign MEM[6841] = MEM[3456] + MEM[3457];
assign MEM[6842] = MEM[3544] + MEM[3545];
assign MEM[6843] = MEM[3687] + MEM[362];
assign MEM[6844] = MEM[3696] + MEM[3697];
assign MEM[6845] = MEM[3711] + MEM[4635];
assign MEM[6846] = MEM[3734] + MEM[1174];
assign MEM[6847] = MEM[3743] + MEM[3079];
assign MEM[6848] = MEM[3776] + MEM[3777];
assign MEM[6849] = MEM[3995] + MEM[4156];
assign MEM[6850] = MEM[4032] + MEM[4033];
assign MEM[6851] = MEM[4034] + MEM[4035];
assign MEM[6852] = MEM[4036] + MEM[6850];
assign MEM[6853] = MEM[4184] + MEM[4185];
assign MEM[6854] = MEM[4208] + MEM[4209];
assign MEM[6855] = MEM[4232] + MEM[4233];
assign MEM[6856] = MEM[4261] + MEM[677];
assign MEM[6857] = MEM[4280] + MEM[4281];
assign MEM[6858] = MEM[4352] + MEM[4353];
assign MEM[6859] = MEM[4424] + MEM[4425];
assign MEM[6860] = MEM[4480] + MEM[4481];
assign MEM[6861] = MEM[4482] + MEM[4483];
assign MEM[6862] = MEM[4484] + MEM[6860];
assign MEM[6863] = MEM[4520] + MEM[4521];
assign MEM[6864] = MEM[4608] + MEM[4609];
assign MEM[6865] = MEM[4688] + MEM[4689];
assign MEM[6866] = MEM[4690] + MEM[6865];
assign MEM[6867] = MEM[4696] + MEM[4697];
assign MEM[6868] = MEM[4698] + MEM[4699];
assign MEM[6869] = MEM[4700] + MEM[6867];
assign MEM[6870] = MEM[4737] + MEM[4736];
assign MEM[6871] = MEM[4776] + MEM[4777];
assign MEM[6872] = MEM[4944] + MEM[4945];
assign MEM[6873] = MEM[5056] + MEM[5058];
assign MEM[6874] = MEM[5096] + MEM[5097];
assign MEM[6875] = MEM[5104] + MEM[5105];
assign MEM[6876] = MEM[5204] + MEM[159];
assign MEM[6877] = MEM[5329] + MEM[5328];
assign MEM[6878] = MEM[5333] + MEM[3052];
assign MEM[6879] = MEM[5336] + MEM[5337];
assign MEM[6880] = MEM[5512] + MEM[5513];
assign MEM[6881] = MEM[5520] + MEM[5521];
assign MEM[6882] = MEM[5608] + MEM[5609];
assign MEM[6883] = MEM[5610] + MEM[5611];
assign MEM[6884] = MEM[5612] + MEM[6882];
assign MEM[6885] = MEM[5672] + MEM[5673];
assign MEM[6886] = MEM[5720] + MEM[5721];
assign MEM[6887] = MEM[5864] + MEM[5865];
assign MEM[6888] = MEM[5920] + MEM[5921];
assign MEM[6889] = MEM[5992] + MEM[5993];
assign MEM[6890] = MEM[6064] + MEM[6065];
assign MEM[6891] = MEM[6066] + MEM[6067];
assign MEM[6892] = MEM[6068] + MEM[6890];
assign MEM[6893] = MEM[6160] + MEM[6161];
assign MEM[6894] = MEM[6208] + MEM[6209];
assign MEM[6895] = MEM[6210] + MEM[6894];
assign MEM[6896] = MEM[6273] + MEM[4756];
assign MEM[6897] = MEM[6275] + MEM[6282];
assign MEM[6898] = MEM[6277] + MEM[6297];
assign MEM[6899] = MEM[6285] + MEM[6294];
assign MEM[6900] = MEM[6757] + MEM[6758];
assign MEM[6901] = MEM[6760] + MEM[6761];
assign MEM[6902] = MEM[6763] + MEM[6764];
assign MEM[6903] = MEM[6766] + MEM[6767];
assign MEM[6904] = MEM[6769] + MEM[6770];
assign MEM[6905] = MEM[6772] + MEM[6773];
assign MEM[6906] = MEM[6781] + MEM[6782];
assign MEM[6907] = MEM[6783] + MEM[482];
assign MEM[6908] = MEM[6789] + MEM[6790];
assign MEM[6909] = MEM[6792] + MEM[6793];
assign MEM[6910] = MEM[6824] + MEM[6825];
assign MEM[6911] = MEM[6830] + MEM[6374];
assign MEM[6912] = MEM[6834] + MEM[6835];
assign MEM[6913] = MEM[6851] + MEM[6852];
assign MEM[6914] = MEM[6861] + MEM[6862];
assign MEM[6915] = MEM[6868] + MEM[6869];
assign MEM[6916] = MEM[6883] + MEM[6884];
assign MEM[6917] = MEM[6891] + MEM[6892];
assign MEM[6918] = MEM[40] + MEM[41];
assign MEM[6919] = MEM[42] + MEM[43];
assign MEM[6920] = MEM[44] + MEM[6918];
assign MEM[6921] = MEM[213] + MEM[5556];
assign MEM[6922] = MEM[300] + MEM[299];
assign MEM[6923] = MEM[355] + MEM[806];
assign MEM[6924] = MEM[414] + MEM[5194];
assign MEM[6925] = MEM[416] + MEM[417];
assign MEM[6926] = MEM[418] + MEM[419];
assign MEM[6927] = MEM[420] + MEM[6925];
assign MEM[6928] = MEM[510] + MEM[626];
assign MEM[6929] = MEM[520] + MEM[521];
assign MEM[6930] = MEM[547] + MEM[3245];
assign MEM[6931] = MEM[560] + MEM[561];
assign MEM[6932] = MEM[624] + MEM[625];
assign MEM[6933] = MEM[632] + MEM[633];
assign MEM[6934] = MEM[664] + MEM[665];
assign MEM[6935] = MEM[666] + MEM[667];
assign MEM[6936] = MEM[668] + MEM[6934];
assign MEM[6937] = MEM[775] + MEM[5263];
assign MEM[6938] = MEM[810] + MEM[2051];
assign MEM[6939] = MEM[1040] + MEM[1041];
assign MEM[6940] = MEM[1152] + MEM[1153];
assign MEM[6941] = MEM[1184] + MEM[1185];
assign MEM[6942] = MEM[1200] + MEM[1201];
assign MEM[6943] = MEM[1232] + MEM[1233];
assign MEM[6944] = MEM[1256] + MEM[1257];
assign MEM[6945] = MEM[1264] + MEM[1265];
assign MEM[6946] = MEM[1304] + MEM[1305];
assign MEM[6947] = MEM[1312] + MEM[1313];
assign MEM[6948] = MEM[1333] + MEM[1189];
assign MEM[6949] = MEM[1341] + MEM[4218];
assign MEM[6950] = MEM[1376] + MEM[1377];
assign MEM[6951] = MEM[1383] + MEM[2955];
assign MEM[6952] = MEM[1448] + MEM[1449];
assign MEM[6953] = MEM[1498] + MEM[6413];
assign MEM[6954] = MEM[1529] + MEM[1528];
assign MEM[6955] = MEM[1536] + MEM[1537];
assign MEM[6956] = MEM[1721] + MEM[1720];
assign MEM[6957] = MEM[1816] + MEM[1817];
assign MEM[6958] = MEM[1825] + MEM[1824];
assign MEM[6959] = MEM[1835] + MEM[2757];
assign MEM[6960] = MEM[1888] + MEM[1889];
assign MEM[6961] = MEM[1910] + MEM[4277];
assign MEM[6962] = MEM[1920] + MEM[1921];
assign MEM[6963] = MEM[1992] + MEM[1993];
assign MEM[6964] = MEM[2048] + MEM[2049];
assign MEM[6965] = MEM[2064] + MEM[2065];
assign MEM[6966] = MEM[2068] + MEM[5279];
assign MEM[6967] = MEM[2094] + MEM[3885];
assign MEM[6968] = MEM[2096] + MEM[2097];
assign MEM[6969] = MEM[2175] + MEM[2748];
assign MEM[6970] = MEM[2201] + MEM[2200];
assign MEM[6971] = MEM[2216] + MEM[2217];
assign MEM[6972] = MEM[2234] + MEM[6664];
assign MEM[6973] = MEM[2305] + MEM[2304];
assign MEM[6974] = MEM[2329] + MEM[2328];
assign MEM[6975] = MEM[2638] + MEM[5573];
assign MEM[6976] = MEM[2639] + MEM[4723];
assign MEM[6977] = MEM[2672] + MEM[2664];
assign MEM[6978] = MEM[2688] + MEM[2689];
assign MEM[6979] = MEM[2690] + MEM[2691];
assign MEM[6980] = MEM[2730] + MEM[3803];
assign MEM[6981] = MEM[2793] + MEM[2792];
assign MEM[6982] = MEM[2832] + MEM[2833];
assign MEM[6983] = MEM[3014] + MEM[1365];
assign MEM[6984] = MEM[3045] + MEM[862];
assign MEM[6985] = MEM[3186] + MEM[3184];
assign MEM[6986] = MEM[3201] + MEM[3200];
assign MEM[6987] = MEM[3291] + MEM[4542];
assign MEM[6988] = MEM[3304] + MEM[3305];
assign MEM[6989] = MEM[3360] + MEM[3361];
assign MEM[6990] = MEM[3362] + MEM[3363];
assign MEM[6991] = MEM[3364] + MEM[6989];
assign MEM[6992] = MEM[3371] + MEM[1895];
assign MEM[6993] = MEM[3402] + MEM[6488];
assign MEM[6994] = MEM[3425] + MEM[3424];
assign MEM[6995] = MEM[3432] + MEM[3433];
assign MEM[6996] = MEM[3454] + MEM[1043];
assign MEM[6997] = MEM[3506] + MEM[6684];
assign MEM[6998] = MEM[3578] + MEM[3004];
assign MEM[6999] = MEM[3720] + MEM[3721];
assign MEM[7000] = MEM[3883] + MEM[3882];
assign MEM[7001] = MEM[3897] + MEM[3896];
assign MEM[7002] = MEM[3912] + MEM[3913];
assign MEM[7003] = MEM[3925] + MEM[2542];
assign MEM[7004] = MEM[3978] + MEM[3954];
assign MEM[7005] = MEM[4016] + MEM[4017];
assign MEM[7006] = MEM[4018] + MEM[515];
assign MEM[7007] = MEM[4024] + MEM[4025];
assign MEM[7008] = MEM[4026] + MEM[4027];
assign MEM[7009] = MEM[4028] + MEM[7007];
assign MEM[7010] = MEM[4056] + MEM[4057];
assign MEM[7011] = MEM[4100] + MEM[2940];
assign MEM[7012] = MEM[4206] + MEM[5893];
assign MEM[7013] = MEM[4254] + MEM[3287];
assign MEM[7014] = MEM[4272] + MEM[4273];
assign MEM[7015] = MEM[4376] + MEM[4377];
assign MEM[7016] = MEM[4440] + MEM[4441];
assign MEM[7017] = MEM[4464] + MEM[4465];
assign MEM[7018] = MEM[4466] + MEM[3213];
assign MEM[7019] = MEM[4488] + MEM[4489];
assign MEM[7020] = MEM[4544] + MEM[4545];
assign MEM[7021] = MEM[4600] + MEM[4602];
assign MEM[7022] = MEM[4720] + MEM[4721];
assign MEM[7023] = MEM[4784] + MEM[4785];
assign MEM[7024] = MEM[4824] + MEM[4825];
assign MEM[7025] = MEM[4830] + MEM[1055];
assign MEM[7026] = MEM[4840] + MEM[4841];
assign MEM[7027] = MEM[4955] + MEM[6123];
assign MEM[7028] = MEM[5057] + MEM[6873];
assign MEM[7029] = MEM[5080] + MEM[5081];
assign MEM[7030] = MEM[5088] + MEM[5089];
assign MEM[7031] = MEM[5176] + MEM[5177];
assign MEM[7032] = MEM[5184] + MEM[5185];
assign MEM[7033] = MEM[5408] + MEM[5409];
assign MEM[7034] = MEM[5433] + MEM[5432];
assign MEM[7035] = MEM[5536] + MEM[5537];
assign MEM[7036] = MEM[5544] + MEM[5545];
assign MEM[7037] = MEM[5568] + MEM[5569];
assign MEM[7038] = MEM[5732] + MEM[6272];
assign MEM[7039] = MEM[5745] + MEM[5744];
assign MEM[7040] = MEM[5822] + MEM[291];
assign MEM[7041] = MEM[5976] + MEM[5977];
assign MEM[7042] = MEM[6124] + MEM[3828];
assign MEM[7043] = MEM[6127] + MEM[85];
assign MEM[7044] = MEM[6144] + MEM[6145];
assign MEM[7045] = MEM[6192] + MEM[6193];
assign MEM[7046] = MEM[6274] + MEM[1075];
assign MEM[7047] = MEM[6281] + MEM[1863];
assign MEM[7048] = MEM[6287] + MEM[6304];
assign MEM[7049] = MEM[6308] + MEM[4925];
assign MEM[7050] = MEM[6312] + MEM[6298];
assign MEM[7051] = MEM[6368] + MEM[2771];
assign MEM[7052] = MEM[6439] + MEM[2035];
assign MEM[7053] = MEM[6919] + MEM[6920];
assign MEM[7054] = MEM[6926] + MEM[6927];
assign MEM[7055] = MEM[6935] + MEM[6936];
assign MEM[7056] = MEM[6978] + MEM[6979];
assign MEM[7057] = MEM[6990] + MEM[6991];
assign MEM[7058] = MEM[7008] + MEM[7009];
assign MEM[7059] = MEM[7010] + MEM[4058];
assign MEM[7060] = MEM[7014] + MEM[4274];
assign MEM[7061] = MEM[7045] + MEM[6194];
assign MEM[7062] = MEM[13] + MEM[1804];
assign MEM[7063] = MEM[276] + MEM[2564];
assign MEM[7064] = MEM[400] + MEM[401];
assign MEM[7065] = MEM[402] + MEM[7064];
assign MEM[7066] = MEM[488] + MEM[489];
assign MEM[7067] = MEM[490] + MEM[491];
assign MEM[7068] = MEM[492] + MEM[7066];
assign MEM[7069] = MEM[589] + MEM[1460];
assign MEM[7070] = MEM[720] + MEM[721];
assign MEM[7071] = MEM[753] + MEM[752];
assign MEM[7072] = MEM[789] + MEM[3407];
assign MEM[7073] = MEM[817] + MEM[816];
assign MEM[7074] = MEM[833] + MEM[832];
assign MEM[7075] = MEM[968] + MEM[969];
assign MEM[7076] = MEM[981] + MEM[1862];
assign MEM[7077] = MEM[1112] + MEM[1113];
assign MEM[7078] = MEM[1114] + MEM[1115];
assign MEM[7079] = MEM[1116] + MEM[7077];
assign MEM[7080] = MEM[1120] + MEM[1121];
assign MEM[7081] = MEM[1122] + MEM[1123];
assign MEM[7082] = MEM[1124] + MEM[7080];
assign MEM[7083] = MEM[1125] + MEM[2428];
assign MEM[7084] = MEM[1210] + MEM[6547];
assign MEM[7085] = MEM[1224] + MEM[1225];
assign MEM[7086] = MEM[1254] + MEM[3555];
assign MEM[7087] = MEM[1328] + MEM[1329];
assign MEM[7088] = MEM[1632] + MEM[1633];
assign MEM[7089] = MEM[1640] + MEM[1641];
assign MEM[7090] = MEM[1676] + MEM[1619];
assign MEM[7091] = MEM[1694] + MEM[1047];
assign MEM[7092] = MEM[1696] + MEM[1697];
assign MEM[7093] = MEM[1856] + MEM[1857];
assign MEM[7094] = MEM[1867] + MEM[1118];
assign MEM[7095] = MEM[1894] + MEM[1421];
assign MEM[7096] = MEM[1928] + MEM[1929];
assign MEM[7097] = MEM[1931] + MEM[1770];
assign MEM[7098] = MEM[1944] + MEM[1945];
assign MEM[7099] = MEM[1961] + MEM[1960];
assign MEM[7100] = MEM[1963] + MEM[2412];
assign MEM[7101] = MEM[1974] + MEM[5902];
assign MEM[7102] = MEM[1979] + MEM[1511];
assign MEM[7103] = MEM[2000] + MEM[2001];
assign MEM[7104] = MEM[2079] + MEM[2644];
assign MEM[7105] = MEM[2133] + MEM[2987];
assign MEM[7106] = MEM[2145] + MEM[2144];
assign MEM[7107] = MEM[2165] + MEM[2670];
assign MEM[7108] = MEM[2176] + MEM[2177];
assign MEM[7109] = MEM[2377] + MEM[2376];
assign MEM[7110] = MEM[2401] + MEM[2400];
assign MEM[7111] = MEM[2433] + MEM[2432];
assign MEM[7112] = MEM[2443] + MEM[1726];
assign MEM[7113] = MEM[2456] + MEM[2457];
assign MEM[7114] = MEM[2458] + MEM[7113];
assign MEM[7115] = MEM[2500] + MEM[1035];
assign MEM[7116] = MEM[2515] + MEM[2587];
assign MEM[7117] = MEM[2521] + MEM[2520];
assign MEM[7118] = MEM[2608] + MEM[2609];
assign MEM[7119] = MEM[2617] + MEM[2616];
assign MEM[7120] = MEM[2625] + MEM[2624];
assign MEM[7121] = MEM[2636] + MEM[3492];
assign MEM[7122] = MEM[2673] + MEM[2674];
assign MEM[7123] = MEM[2685] + MEM[3562];
assign MEM[7124] = MEM[2805] + MEM[999];
assign MEM[7125] = MEM[2824] + MEM[2825];
assign MEM[7126] = MEM[2911] + MEM[4299];
assign MEM[7127] = MEM[2992] + MEM[2993];
assign MEM[7128] = MEM[3017] + MEM[3016];
assign MEM[7129] = MEM[3050] + MEM[6829];
assign MEM[7130] = MEM[3191] + MEM[2374];
assign MEM[7131] = MEM[3376] + MEM[3377];
assign MEM[7132] = MEM[3378] + MEM[7131];
assign MEM[7133] = MEM[3386] + MEM[1755];
assign MEM[7134] = MEM[3568] + MEM[3569];
assign MEM[7135] = MEM[3664] + MEM[3665];
assign MEM[7136] = MEM[3673] + MEM[3672];
assign MEM[7137] = MEM[3682] + MEM[46];
assign MEM[7138] = MEM[3712] + MEM[3713];
assign MEM[7139] = MEM[3738] + MEM[3962];
assign MEM[7140] = MEM[3768] + MEM[3769];
assign MEM[7141] = MEM[3784] + MEM[3785];
assign MEM[7142] = MEM[3798] + MEM[4644];
assign MEM[7143] = MEM[3831] + MEM[1655];
assign MEM[7144] = MEM[4106] + MEM[4107];
assign MEM[7145] = MEM[4114] + MEM[6069];
assign MEM[7146] = MEM[4117] + MEM[3206];
assign MEM[7147] = MEM[4144] + MEM[4145];
assign MEM[7148] = MEM[4192] + MEM[4193];
assign MEM[7149] = MEM[4228] + MEM[108];
assign MEM[7150] = MEM[4368] + MEM[4369];
assign MEM[7151] = MEM[4378] + MEM[7015];
assign MEM[7152] = MEM[4601] + MEM[7021];
assign MEM[7153] = MEM[4623] + MEM[102];
assign MEM[7154] = MEM[4651] + MEM[4349];
assign MEM[7155] = MEM[4680] + MEM[4681];
assign MEM[7156] = MEM[4704] + MEM[4705];
assign MEM[7157] = MEM[4706] + MEM[4707];
assign MEM[7158] = MEM[4708] + MEM[7156];
assign MEM[7159] = MEM[4709] + MEM[590];
assign MEM[7160] = MEM[4792] + MEM[4793];
assign MEM[7161] = MEM[4947] + MEM[5723];
assign MEM[7162] = MEM[4971] + MEM[523];
assign MEM[7163] = MEM[5000] + MEM[5001];
assign MEM[7164] = MEM[5024] + MEM[5025];
assign MEM[7165] = MEM[5128] + MEM[5129];
assign MEM[7166] = MEM[5178] + MEM[797];
assign MEM[7167] = MEM[5357] + MEM[4372];
assign MEM[7168] = MEM[5464] + MEM[5465];
assign MEM[7169] = MEM[5505] + MEM[5504];
assign MEM[7170] = MEM[5532] + MEM[3932];
assign MEM[7171] = MEM[5554] + MEM[4387];
assign MEM[7172] = MEM[5560] + MEM[5561];
assign MEM[7173] = MEM[5572] + MEM[1787];
assign MEM[7174] = MEM[5624] + MEM[5625];
assign MEM[7175] = MEM[5626] + MEM[7174];
assign MEM[7176] = MEM[5664] + MEM[5665];
assign MEM[7177] = MEM[5688] + MEM[5689];
assign MEM[7178] = MEM[5729] + MEM[5728];
assign MEM[7179] = MEM[5758] + MEM[3773];
assign MEM[7180] = MEM[5781] + MEM[5327];
assign MEM[7181] = MEM[5808] + MEM[5809];
assign MEM[7182] = MEM[5810] + MEM[5811];
assign MEM[7183] = MEM[5812] + MEM[7181];
assign MEM[7184] = MEM[5896] + MEM[6283];
assign MEM[7185] = MEM[6040] + MEM[6041];
assign MEM[7186] = MEM[6042] + MEM[6043];
assign MEM[7187] = MEM[6044] + MEM[7185];
assign MEM[7188] = MEM[6056] + MEM[6057];
assign MEM[7189] = MEM[6058] + MEM[6059];
assign MEM[7190] = MEM[6060] + MEM[7188];
assign MEM[7191] = MEM[6183] + MEM[2708];
assign MEM[7192] = MEM[6184] + MEM[6185];
assign MEM[7193] = MEM[6238] + MEM[636];
assign MEM[7194] = MEM[6256] + MEM[6257];
assign MEM[7195] = MEM[6258] + MEM[6259];
assign MEM[7196] = MEM[6260] + MEM[7194];
assign MEM[7197] = MEM[6279] + MEM[205];
assign MEM[7198] = MEM[6286] + MEM[3986];
assign MEM[7199] = MEM[6289] + MEM[4135];
assign MEM[7200] = MEM[6293] + MEM[5805];
assign MEM[7201] = MEM[6299] + MEM[5198];
assign MEM[7202] = MEM[6302] + MEM[6338];
assign MEM[7203] = MEM[6322] + MEM[6353];
assign MEM[7204] = MEM[6331] + MEM[2619];
assign MEM[7205] = MEM[6344] + MEM[2854];
assign MEM[7206] = MEM[6363] + MEM[2346];
assign MEM[7207] = MEM[7067] + MEM[7068];
assign MEM[7208] = MEM[7078] + MEM[7079];
assign MEM[7209] = MEM[7081] + MEM[7082];
assign MEM[7210] = MEM[7136] + MEM[3674];
assign MEM[7211] = MEM[7157] + MEM[7158];
assign MEM[7212] = MEM[7163] + MEM[5002];
assign MEM[7213] = MEM[7164] + MEM[5026];
assign MEM[7214] = MEM[7168] + MEM[5466];
assign MEM[7215] = MEM[7182] + MEM[7183];
assign MEM[7216] = MEM[7186] + MEM[7187];
assign MEM[7217] = MEM[7189] + MEM[7190];
assign MEM[7218] = MEM[7195] + MEM[7196];
assign MEM[7219] = MEM[6] + MEM[3005];
assign MEM[7220] = MEM[56] + MEM[57];
assign MEM[7221] = MEM[58] + MEM[59];
assign MEM[7222] = MEM[60] + MEM[7220];
assign MEM[7223] = MEM[104] + MEM[105];
assign MEM[7224] = MEM[106] + MEM[7223];
assign MEM[7225] = MEM[181] + MEM[535];
assign MEM[7226] = MEM[184] + MEM[185];
assign MEM[7227] = MEM[186] + MEM[187];
assign MEM[7228] = MEM[188] + MEM[7226];
assign MEM[7229] = MEM[208] + MEM[209];
assign MEM[7230] = MEM[210] + MEM[211];
assign MEM[7231] = MEM[212] + MEM[7229];
assign MEM[7232] = MEM[312] + MEM[313];
assign MEM[7233] = MEM[376] + MEM[377];
assign MEM[7234] = MEM[446] + MEM[932];
assign MEM[7235] = MEM[494] + MEM[558];
assign MEM[7236] = MEM[614] + MEM[1387];
assign MEM[7237] = MEM[616] + MEM[617];
assign MEM[7238] = MEM[643] + MEM[2211];
assign MEM[7239] = MEM[719] + MEM[175];
assign MEM[7240] = MEM[874] + MEM[1999];
assign MEM[7241] = MEM[901] + MEM[917];
assign MEM[7242] = MEM[902] + MEM[2724];
assign MEM[7243] = MEM[1074] + MEM[3844];
assign MEM[7244] = MEM[1134] + MEM[1037];
assign MEM[7245] = MEM[1159] + MEM[980];
assign MEM[7246] = MEM[1243] + MEM[1638];
assign MEM[7247] = MEM[1301] + MEM[1518];
assign MEM[7248] = MEM[1324] + MEM[2804];
assign MEM[7249] = MEM[1471] + MEM[2613];
assign MEM[7250] = MEM[1552] + MEM[1553];
assign MEM[7251] = MEM[1560] + MEM[1561];
assign MEM[7252] = MEM[1562] + MEM[7251];
assign MEM[7253] = MEM[1584] + MEM[1585];
assign MEM[7254] = MEM[1586] + MEM[7253];
assign MEM[7255] = MEM[1600] + MEM[1601];
assign MEM[7256] = MEM[1604] + MEM[110];
assign MEM[7257] = MEM[1652] + MEM[3791];
assign MEM[7258] = MEM[1688] + MEM[1689];
assign MEM[7259] = MEM[1712] + MEM[1713];
assign MEM[7260] = MEM[1797] + MEM[1829];
assign MEM[7261] = MEM[1896] + MEM[1897];
assign MEM[7262] = MEM[1912] + MEM[1913];
assign MEM[7263] = MEM[2016] + MEM[2017];
assign MEM[7264] = MEM[2018] + MEM[2019];
assign MEM[7265] = MEM[2020] + MEM[7263];
assign MEM[7266] = MEM[2024] + MEM[2025];
assign MEM[7267] = MEM[2026] + MEM[2027];
assign MEM[7268] = MEM[2085] + MEM[3618];
assign MEM[7269] = MEM[2138] + MEM[4381];
assign MEM[7270] = MEM[2141] + MEM[4219];
assign MEM[7271] = MEM[2151] + MEM[2997];
assign MEM[7272] = MEM[2209] + MEM[2208];
assign MEM[7273] = MEM[2272] + MEM[2273];
assign MEM[7274] = MEM[2288] + MEM[2289];
assign MEM[7275] = MEM[2482] + MEM[4619];
assign MEM[7276] = MEM[2562] + MEM[1407];
assign MEM[7277] = MEM[2600] + MEM[2601];
assign MEM[7278] = MEM[2642] + MEM[6366];
assign MEM[7279] = MEM[2719] + MEM[2055];
assign MEM[7280] = MEM[2777] + MEM[2776];
assign MEM[7281] = MEM[2818] + MEM[109];
assign MEM[7282] = MEM[2848] + MEM[2849];
assign MEM[7283] = MEM[2978] + MEM[3970];
assign MEM[7284] = MEM[3024] + MEM[3025];
assign MEM[7285] = MEM[3033] + MEM[3032];
assign MEM[7286] = MEM[3066] + MEM[5323];
assign MEM[7287] = MEM[3240] + MEM[3241];
assign MEM[7288] = MEM[3248] + MEM[3249];
assign MEM[7289] = MEM[3255] + MEM[3949];
assign MEM[7290] = MEM[3256] + MEM[3258];
assign MEM[7291] = MEM[3389] + MEM[5061];
assign MEM[7292] = MEM[3406] + MEM[4811];
assign MEM[7293] = MEM[3430] + MEM[4674];
assign MEM[7294] = MEM[3455] + MEM[3612];
assign MEM[7295] = MEM[3531] + MEM[4103];
assign MEM[7296] = MEM[3635] + MEM[2421];
assign MEM[7297] = MEM[3637] + MEM[381];
assign MEM[7298] = MEM[3707] + MEM[5443];
assign MEM[7299] = MEM[3730] + MEM[3498];
assign MEM[7300] = MEM[3732] + MEM[3316];
assign MEM[7301] = MEM[3750] + MEM[1956];
assign MEM[7302] = MEM[3760] + MEM[3761];
assign MEM[7303] = MEM[3824] + MEM[3825];
assign MEM[7304] = MEM[3876] + MEM[4603];
assign MEM[7305] = MEM[3887] + MEM[1691];
assign MEM[7306] = MEM[3947] + MEM[5205];
assign MEM[7307] = MEM[3982] + MEM[686];
assign MEM[7308] = MEM[3988] + MEM[2302];
assign MEM[7309] = MEM[4160] + MEM[4161];
assign MEM[7310] = MEM[4171] + MEM[3070];
assign MEM[7311] = MEM[4198] + MEM[755];
assign MEM[7312] = MEM[4240] + MEM[4241];
assign MEM[7313] = MEM[4298] + MEM[4583];
assign MEM[7314] = MEM[4300] + MEM[5483];
assign MEM[7315] = MEM[4325] + MEM[631];
assign MEM[7316] = MEM[4383] + MEM[292];
assign MEM[7317] = MEM[4404] + MEM[3767];
assign MEM[7318] = MEM[4446] + MEM[4683];
assign MEM[7319] = MEM[4616] + MEM[4617];
assign MEM[7320] = MEM[4643] + MEM[3365];
assign MEM[7321] = MEM[4758] + MEM[4755];
assign MEM[7322] = MEM[4797] + MEM[4397];
assign MEM[7323] = MEM[4800] + MEM[4801];
assign MEM[7324] = MEM[4812] + MEM[5685];
assign MEM[7325] = MEM[4880] + MEM[4881];
assign MEM[7326] = MEM[4981] + MEM[539];
assign MEM[7327] = MEM[4984] + MEM[4985];
assign MEM[7328] = MEM[4992] + MEM[4993];
assign MEM[7329] = MEM[4996] + MEM[3495];
assign MEM[7330] = MEM[5036] + MEM[335];
assign MEM[7331] = MEM[5064] + MEM[5065];
assign MEM[7332] = MEM[5130] + MEM[7165];
assign MEM[7333] = MEM[5224] + MEM[5225];
assign MEM[7334] = MEM[5264] + MEM[5265];
assign MEM[7335] = MEM[5268] + MEM[1220];
assign MEM[7336] = MEM[5272] + MEM[5273];
assign MEM[7337] = MEM[5311] + MEM[502];
assign MEM[7338] = MEM[5319] + MEM[3748];
assign MEM[7339] = MEM[5400] + MEM[5401];
assign MEM[7340] = MEM[5441] + MEM[5440];
assign MEM[7341] = MEM[5480] + MEM[5481];
assign MEM[7342] = MEM[5488] + MEM[5489];
assign MEM[7343] = MEM[5510] + MEM[2949];
assign MEM[7344] = MEM[5606] + MEM[1171];
assign MEM[7345] = MEM[5607] + MEM[1540];
assign MEM[7346] = MEM[5616] + MEM[5617];
assign MEM[7347] = MEM[5618] + MEM[5619];
assign MEM[7348] = MEM[5620] + MEM[7346];
assign MEM[7349] = MEM[5648] + MEM[5649];
assign MEM[7350] = MEM[5807] + MEM[5418];
assign MEM[7351] = MEM[5871] + MEM[1871];
assign MEM[7352] = MEM[5897] + MEM[6325];
assign MEM[7353] = MEM[5899] + MEM[1086];
assign MEM[7354] = MEM[5916] + MEM[3325];
assign MEM[7355] = MEM[5926] + MEM[2014];
assign MEM[7356] = MEM[5969] + MEM[5968];
assign MEM[7357] = MEM[5982] + MEM[559];
assign MEM[7358] = MEM[5984] + MEM[5985];
assign MEM[7359] = MEM[5990] + MEM[2501];
assign MEM[7360] = MEM[6032] + MEM[6033];
assign MEM[7361] = MEM[6034] + MEM[6035];
assign MEM[7362] = MEM[6036] + MEM[7360];
assign MEM[7363] = MEM[6136] + MEM[6137];
assign MEM[7364] = MEM[6146] + MEM[7044];
assign MEM[7365] = MEM[6176] + MEM[6177];
assign MEM[7366] = MEM[6186] + MEM[7192];
assign MEM[7367] = MEM[6261] + MEM[4847];
assign MEM[7368] = MEM[6290] + MEM[2939];
assign MEM[7369] = MEM[6291] + MEM[909];
assign MEM[7370] = MEM[6295] + MEM[4270];
assign MEM[7371] = MEM[6296] + MEM[3244];
assign MEM[7372] = MEM[6300] + MEM[1261];
assign MEM[7373] = MEM[6301] + MEM[735];
assign MEM[7374] = MEM[6309] + MEM[4074];
assign MEM[7375] = MEM[6311] + MEM[5838];
assign MEM[7376] = MEM[6317] + MEM[4974];
assign MEM[7377] = MEM[6333] + MEM[4694];
assign MEM[7378] = MEM[6337] + MEM[5986];
assign MEM[7379] = MEM[6339] + MEM[6340];
assign MEM[7380] = MEM[6345] + MEM[2882];
assign MEM[7381] = MEM[6364] + MEM[780];
assign MEM[7382] = MEM[6369] + MEM[6328];
assign MEM[7383] = MEM[6373] + MEM[2979];
assign MEM[7384] = MEM[6375] + MEM[3322];
assign MEM[7385] = MEM[6453] + MEM[6303];
assign MEM[7386] = MEM[7221] + MEM[7222];
assign MEM[7387] = MEM[7227] + MEM[7228];
assign MEM[7388] = MEM[7230] + MEM[7231];
assign MEM[7389] = MEM[7232] + MEM[314];
assign MEM[7390] = MEM[7264] + MEM[7265];
assign MEM[7391] = MEM[7266] + MEM[7267];
assign MEM[7392] = MEM[7309] + MEM[4162];
assign MEM[7393] = MEM[7313] + MEM[6315];
assign MEM[7394] = MEM[7347] + MEM[7348];
assign MEM[7395] = MEM[7361] + MEM[7362];
assign MEM[7396] = MEM[24] + MEM[25];
assign MEM[7397] = MEM[26] + MEM[27];
assign MEM[7398] = MEM[28] + MEM[7396];
assign MEM[7399] = MEM[78] + MEM[5861];
assign MEM[7400] = MEM[80] + MEM[81];
assign MEM[7401] = MEM[82] + MEM[83];
assign MEM[7402] = MEM[84] + MEM[7400];
assign MEM[7403] = MEM[189] + MEM[3630];
assign MEM[7404] = MEM[240] + MEM[241];
assign MEM[7405] = MEM[242] + MEM[243];
assign MEM[7406] = MEM[244] + MEM[7404];
assign MEM[7407] = MEM[254] + MEM[3655];
assign MEM[7408] = MEM[280] + MEM[281];
assign MEM[7409] = MEM[282] + MEM[7408];
assign MEM[7410] = MEM[287] + MEM[661];
assign MEM[7411] = MEM[347] + MEM[2798];
assign MEM[7412] = MEM[408] + MEM[409];
assign MEM[7413] = MEM[410] + MEM[7412];
assign MEM[7414] = MEM[422] + MEM[2404];
assign MEM[7415] = MEM[448] + MEM[449];
assign MEM[7416] = MEM[450] + MEM[451];
assign MEM[7417] = MEM[452] + MEM[7415];
assign MEM[7418] = MEM[499] + MEM[1700];
assign MEM[7419] = MEM[525] + MEM[4006];
assign MEM[7420] = MEM[566] + MEM[2419];
assign MEM[7421] = MEM[573] + MEM[1502];
assign MEM[7422] = MEM[592] + MEM[593];
assign MEM[7423] = MEM[605] + MEM[3718];
assign MEM[7424] = MEM[635] + MEM[870];
assign MEM[7425] = MEM[688] + MEM[689];
assign MEM[7426] = MEM[690] + MEM[691];
assign MEM[7427] = MEM[692] + MEM[7425];
assign MEM[7428] = MEM[711] + MEM[1765];
assign MEM[7429] = MEM[716] + MEM[926];
assign MEM[7430] = MEM[723] + MEM[3246];
assign MEM[7431] = MEM[734] + MEM[1051];
assign MEM[7432] = MEM[767] + MEM[461];
assign MEM[7433] = MEM[795] + MEM[4975];
assign MEM[7434] = MEM[1008] + MEM[1009];
assign MEM[7435] = MEM[1048] + MEM[1049];
assign MEM[7436] = MEM[1058] + MEM[3029];
assign MEM[7437] = MEM[1104] + MEM[1105];
assign MEM[7438] = MEM[1165] + MEM[565];
assign MEM[7439] = MEM[1194] + MEM[6800];
assign MEM[7440] = MEM[1212] + MEM[779];
assign MEM[7441] = MEM[1213] + MEM[3387];
assign MEM[7442] = MEM[1244] + MEM[3067];
assign MEM[7443] = MEM[1330] + MEM[6334];
assign MEM[7444] = MEM[1368] + MEM[1369];
assign MEM[7445] = MEM[1427] + MEM[5074];
assign MEM[7446] = MEM[1432] + MEM[1433];
assign MEM[7447] = MEM[1443] + MEM[1442];
assign MEM[7448] = MEM[1557] + MEM[1951];
assign MEM[7449] = MEM[1680] + MEM[1681];
assign MEM[7450] = MEM[1695] + MEM[198];
assign MEM[7451] = MEM[1698] + MEM[7092];
assign MEM[7452] = MEM[1704] + MEM[1705];
assign MEM[7453] = MEM[1709] + MEM[5283];
assign MEM[7454] = MEM[1730] + MEM[2765];
assign MEM[7455] = MEM[1772] + MEM[1748];
assign MEM[7456] = MEM[1779] + MEM[437];
assign MEM[7457] = MEM[1814] + MEM[1943];
assign MEM[7458] = MEM[1822] + MEM[2700];
assign MEM[7459] = MEM[1848] + MEM[1849];
assign MEM[7460] = MEM[1858] + MEM[7093];
assign MEM[7461] = MEM[1908] + MEM[3919];
assign MEM[7462] = MEM[1954] + MEM[6318];
assign MEM[7463] = MEM[1964] + MEM[4757];
assign MEM[7464] = MEM[1972] + MEM[3987];
assign MEM[7465] = MEM[1985] + MEM[1984];
assign MEM[7466] = MEM[2008] + MEM[2009];
assign MEM[7467] = MEM[2010] + MEM[7466];
assign MEM[7468] = MEM[2042] + MEM[5171];
assign MEM[7469] = MEM[2066] + MEM[6965];
assign MEM[7470] = MEM[2072] + MEM[2073];
assign MEM[7471] = MEM[2081] + MEM[2080];
assign MEM[7472] = MEM[2221] + MEM[1038];
assign MEM[7473] = MEM[2240] + MEM[2241];
assign MEM[7474] = MEM[2242] + MEM[2243];
assign MEM[7475] = MEM[2244] + MEM[7473];
assign MEM[7476] = MEM[2264] + MEM[2265];
assign MEM[7477] = MEM[2296] + MEM[2297];
assign MEM[7478] = MEM[2319] + MEM[5079];
assign MEM[7479] = MEM[2429] + MEM[1919];
assign MEM[7480] = MEM[2448] + MEM[2449];
assign MEM[7481] = MEM[2503] + MEM[2675];
assign MEM[7482] = MEM[2518] + MEM[4550];
assign MEM[7483] = MEM[2538] + MEM[2546];
assign MEM[7484] = MEM[2563] + MEM[2591];
assign MEM[7485] = MEM[2579] + MEM[1811];
assign MEM[7486] = MEM[2656] + MEM[2665];
assign MEM[7487] = MEM[2680] + MEM[2681];
assign MEM[7488] = MEM[2682] + MEM[2683];
assign MEM[7489] = MEM[2746] + MEM[6332];
assign MEM[7490] = MEM[2770] + MEM[1366];
assign MEM[7491] = MEM[2863] + MEM[2311];
assign MEM[7492] = MEM[2912] + MEM[2913];
assign MEM[7493] = MEM[2914] + MEM[2915];
assign MEM[7494] = MEM[2916] + MEM[7492];
assign MEM[7495] = MEM[2919] + MEM[3314];
assign MEM[7496] = MEM[3002] + MEM[6676];
assign MEM[7497] = MEM[3041] + MEM[3040];
assign MEM[7498] = MEM[3063] + MEM[4284];
assign MEM[7499] = MEM[3142] + MEM[3514];
assign MEM[7500] = MEM[3207] + MEM[310];
assign MEM[7501] = MEM[3211] + MEM[1478];
assign MEM[7502] = MEM[3216] + MEM[3217];
assign MEM[7503] = MEM[3257] + MEM[7290];
assign MEM[7504] = MEM[3338] + MEM[5479];
assign MEM[7505] = MEM[3464] + MEM[3465];
assign MEM[7506] = MEM[3480] + MEM[3481];
assign MEM[7507] = MEM[3574] + MEM[4116];
assign MEM[7508] = MEM[3600] + MEM[3601];
assign MEM[7509] = MEM[3629] + MEM[4692];
assign MEM[7510] = MEM[3688] + MEM[3689];
assign MEM[7511] = MEM[3746] + MEM[6306];
assign MEM[7512] = MEM[3797] + MEM[2339];
assign MEM[7513] = MEM[3808] + MEM[3809];
assign MEM[7514] = MEM[3810] + MEM[3811];
assign MEM[7515] = MEM[3812] + MEM[7513];
assign MEM[7516] = MEM[3890] + MEM[811];
assign MEM[7517] = MEM[3958] + MEM[1447];
assign MEM[7518] = MEM[3981] + MEM[4045];
assign MEM[7519] = MEM[4002] + MEM[3526];
assign MEM[7520] = MEM[4038] + MEM[4746];
assign MEM[7521] = MEM[4048] + MEM[4049];
assign MEM[7522] = MEM[4090] + MEM[6313];
assign MEM[7523] = MEM[4098] + MEM[6005];
assign MEM[7524] = MEM[4234] + MEM[4242];
assign MEM[7525] = MEM[4256] + MEM[4257];
assign MEM[7526] = MEM[4258] + MEM[4259];
assign MEM[7527] = MEM[4260] + MEM[7525];
assign MEM[7528] = MEM[4285] + MEM[3597];
assign MEM[7529] = MEM[4306] + MEM[4307];
assign MEM[7530] = MEM[4360] + MEM[4361];
assign MEM[7531] = MEM[4370] + MEM[7150];
assign MEM[7532] = MEM[4374] + MEM[2348];
assign MEM[7533] = MEM[4392] + MEM[4393];
assign MEM[7534] = MEM[4400] + MEM[4401];
assign MEM[7535] = MEM[4453] + MEM[253];
assign MEM[7536] = MEM[4456] + MEM[4457];
assign MEM[7537] = MEM[4485] + MEM[637];
assign MEM[7538] = MEM[4524] + MEM[479];
assign MEM[7539] = MEM[4554] + MEM[6704];
assign MEM[7540] = MEM[4556] + MEM[1789];
assign MEM[7541] = MEM[4558] + MEM[1693];
assign MEM[7542] = MEM[4584] + MEM[4586];
assign MEM[7543] = MEM[4592] + MEM[4594];
assign MEM[7544] = MEM[4611] + MEM[4610];
assign MEM[7545] = MEM[4622] + MEM[5375];
assign MEM[7546] = MEM[4668] + MEM[1083];
assign MEM[7547] = MEM[4747] + MEM[4883];
assign MEM[7548] = MEM[4768] + MEM[4769];
assign MEM[7549] = MEM[4788] + MEM[1379];
assign MEM[7550] = MEM[4823] + MEM[5179];
assign MEM[7551] = MEM[4888] + MEM[4889];
assign MEM[7552] = MEM[4896] + MEM[4897];
assign MEM[7553] = MEM[4928] + MEM[4929];
assign MEM[7554] = MEM[4930] + MEM[4931];
assign MEM[7555] = MEM[4932] + MEM[7553];
assign MEM[7556] = MEM[4936] + MEM[4937];
assign MEM[7557] = MEM[4938] + MEM[4939];
assign MEM[7558] = MEM[4940] + MEM[7556];
assign MEM[7559] = MEM[4941] + MEM[4230];
assign MEM[7560] = MEM[4952] + MEM[4953];
assign MEM[7561] = MEM[5048] + MEM[5049];
assign MEM[7562] = MEM[5063] + MEM[2972];
assign MEM[7563] = MEM[5152] + MEM[5153];
assign MEM[7564] = MEM[5154] + MEM[5155];
assign MEM[7565] = MEM[5156] + MEM[7563];
assign MEM[7566] = MEM[5281] + MEM[5280];
assign MEM[7567] = MEM[5344] + MEM[5345];
assign MEM[7568] = MEM[5367] + MEM[2758];
assign MEM[7569] = MEM[5419] + MEM[1299];
assign MEM[7570] = MEM[5448] + MEM[5449];
assign MEM[7571] = MEM[5456] + MEM[5457];
assign MEM[7572] = MEM[5482] + MEM[7341];
assign MEM[7573] = MEM[5490] + MEM[7342];
assign MEM[7574] = MEM[5555] + MEM[4492];
assign MEM[7575] = MEM[5576] + MEM[5577];
assign MEM[7576] = MEM[5578] + MEM[7575];
assign MEM[7577] = MEM[5582] + MEM[5638];
assign MEM[7578] = MEM[5656] + MEM[5657];
assign MEM[7579] = MEM[5663] + MEM[1278];
assign MEM[7580] = MEM[5671] + MEM[4679];
assign MEM[7581] = MEM[5741] + MEM[3013];
assign MEM[7582] = MEM[5792] + MEM[5793];
assign MEM[7583] = MEM[5824] + MEM[5825];
assign MEM[7584] = MEM[5826] + MEM[5827];
assign MEM[7585] = MEM[5828] + MEM[7583];
assign MEM[7586] = MEM[5848] + MEM[5849];
assign MEM[7587] = MEM[5850] + MEM[5851];
assign MEM[7588] = MEM[5852] + MEM[7586];
assign MEM[7589] = MEM[5862] + MEM[5947];
assign MEM[7590] = MEM[5994] + MEM[1532];
assign MEM[7591] = MEM[6112] + MEM[6113];
assign MEM[7592] = MEM[6114] + MEM[7591];
assign MEM[7593] = MEM[6132] + MEM[3173];
assign MEM[7594] = MEM[6288] + MEM[2486];
assign MEM[7595] = MEM[6307] + MEM[3090];
assign MEM[7596] = MEM[6310] + MEM[6428];
assign MEM[7597] = MEM[6323] + MEM[2398];
assign MEM[7598] = MEM[6335] + MEM[2111];
assign MEM[7599] = MEM[6341] + MEM[2300];
assign MEM[7600] = MEM[6346] + MEM[6597];
assign MEM[7601] = MEM[6347] + MEM[3290];
assign MEM[7602] = MEM[6359] + MEM[1207];
assign MEM[7603] = MEM[6362] + MEM[6410];
assign MEM[7604] = MEM[6367] + MEM[2747];
assign MEM[7605] = MEM[6370] + MEM[3813];
assign MEM[7606] = MEM[6372] + MEM[2917];
assign MEM[7607] = MEM[6377] + MEM[5891];
assign MEM[7608] = MEM[6381] + MEM[5211];
assign MEM[7609] = MEM[6425] + MEM[3867];
assign MEM[7610] = MEM[6821] + MEM[2554];
assign MEM[7611] = MEM[7135] + MEM[3666];
assign MEM[7612] = MEM[7363] + MEM[6138];
assign MEM[7613] = MEM[7397] + MEM[7398];
assign MEM[7614] = MEM[7401] + MEM[7402];
assign MEM[7615] = MEM[7405] + MEM[7406];
assign MEM[7616] = MEM[7416] + MEM[7417];
assign MEM[7617] = MEM[7426] + MEM[7427];
assign MEM[7618] = MEM[7437] + MEM[1106];
assign MEM[7619] = MEM[7444] + MEM[1370];
assign MEM[7620] = MEM[7447] + MEM[6467];
assign MEM[7621] = MEM[7474] + MEM[7475];
assign MEM[7622] = MEM[7487] + MEM[7488];
assign MEM[7623] = MEM[7493] + MEM[7494];
assign MEM[7624] = MEM[7514] + MEM[7515];
assign MEM[7625] = MEM[7521] + MEM[4050];
assign MEM[7626] = MEM[7526] + MEM[7527];
assign MEM[7627] = MEM[7544] + MEM[6864];
assign MEM[7628] = MEM[7554] + MEM[7555];
assign MEM[7629] = MEM[7557] + MEM[7558];
assign MEM[7630] = MEM[7564] + MEM[7565];
assign MEM[7631] = MEM[7582] + MEM[5794];
assign MEM[7632] = MEM[7584] + MEM[7585];
assign MEM[7633] = MEM[7587] + MEM[7588];
assign MEM[7634] = MEM[0] + MEM[1];
assign MEM[7635] = MEM[2] + MEM[3];
assign MEM[7636] = MEM[4] + MEM[7634];
assign MEM[7637] = MEM[16] + MEM[17];
assign MEM[7638] = MEM[18] + MEM[19];
assign MEM[7639] = MEM[20] + MEM[7637];
assign MEM[7640] = MEM[32] + MEM[33];
assign MEM[7641] = MEM[34] + MEM[35];
assign MEM[7642] = MEM[36] + MEM[7640];
assign MEM[7643] = MEM[37] + MEM[2362];
assign MEM[7644] = MEM[61] + MEM[4667];
assign MEM[7645] = MEM[141] + MEM[4642];
assign MEM[7646] = MEM[229] + MEM[2106];
assign MEM[7647] = MEM[270] + MEM[6045];
assign MEM[7648] = MEM[333] + MEM[4059];
assign MEM[7649] = MEM[365] + MEM[550];
assign MEM[7650] = MEM[370] + MEM[1661];
assign MEM[7651] = MEM[438] + MEM[651];
assign MEM[7652] = MEM[445] + MEM[1229];
assign MEM[7653] = MEM[487] + MEM[1373];
assign MEM[7654] = MEM[514] + MEM[1499];
assign MEM[7655] = MEM[517] + MEM[2635];
assign MEM[7656] = MEM[530] + MEM[2628];
assign MEM[7657] = MEM[531] + MEM[2548];
assign MEM[7658] = MEM[534] + MEM[1639];
assign MEM[7659] = MEM[555] + MEM[2678];
assign MEM[7660] = MEM[581] + MEM[5502];
assign MEM[7661] = MEM[608] + MEM[609];
assign MEM[7662] = MEM[615] + MEM[4551];
assign MEM[7663] = MEM[693] + MEM[1614];
assign MEM[7664] = MEM[702] + MEM[1420];
assign MEM[7665] = MEM[704] + MEM[705];
assign MEM[7666] = MEM[706] + MEM[707];
assign MEM[7667] = MEM[708] + MEM[7665];
assign MEM[7668] = MEM[801] + MEM[800];
assign MEM[7669] = MEM[812] + MEM[4350];
assign MEM[7670] = MEM[827] + MEM[5077];
assign MEM[7671] = MEM[863] + MEM[852];
assign MEM[7672] = MEM[864] + MEM[865];
assign MEM[7673] = MEM[877] + MEM[6348];
assign MEM[7674] = MEM[925] + MEM[1854];
assign MEM[7675] = MEM[946] + MEM[1391];
assign MEM[7676] = MEM[1004] + MEM[2498];
assign MEM[7677] = MEM[1017] + MEM[1016];
assign MEM[7678] = MEM[1163] + MEM[4066];
assign MEM[7679] = MEM[1216] + MEM[1217];
assign MEM[7680] = MEM[1248] + MEM[1249];
assign MEM[7681] = MEM[1252] + MEM[3549];
assign MEM[7682] = MEM[1272] + MEM[1273];
assign MEM[7683] = MEM[1290] + MEM[543];
assign MEM[7684] = MEM[1291] + MEM[2699];
assign MEM[7685] = MEM[1316] + MEM[2654];
assign MEM[7686] = MEM[1343] + MEM[4093];
assign MEM[7687] = MEM[1381] + MEM[3303];
assign MEM[7688] = MEM[1431] + MEM[1463];
assign MEM[7689] = MEM[1452] + MEM[1103];
assign MEM[7690] = MEM[1472] + MEM[1473];
assign MEM[7691] = MEM[1480] + MEM[1481];
assign MEM[7692] = MEM[1491] + MEM[5708];
assign MEM[7693] = MEM[1492] + MEM[1847];
assign MEM[7694] = MEM[1630] + MEM[1916];
assign MEM[7695] = MEM[1636] + MEM[4463];
assign MEM[7696] = MEM[1664] + MEM[1665];
assign MEM[7697] = MEM[1675] + MEM[1674];
assign MEM[7698] = MEM[1686] + MEM[3132];
assign MEM[7699] = MEM[1737] + MEM[1736];
assign MEM[7700] = MEM[1767] + MEM[3292];
assign MEM[7701] = MEM[1776] + MEM[1777];
assign MEM[7702] = MEM[1781] + MEM[2195];
assign MEM[7703] = MEM[1791] + MEM[6157];
assign MEM[7704] = MEM[1805] + MEM[1739];
assign MEM[7705] = MEM[1851] + MEM[3647];
assign MEM[7706] = MEM[1880] + MEM[1881];
assign MEM[7707] = MEM[1893] + MEM[4231];
assign MEM[7708] = MEM[1904] + MEM[1905];
assign MEM[7709] = MEM[1973] + MEM[4566];
assign MEM[7710] = MEM[2011] + MEM[2357];
assign MEM[7711] = MEM[2034] + MEM[6148];
assign MEM[7712] = MEM[2060] + MEM[5350];
assign MEM[7713] = MEM[2143] + MEM[5099];
assign MEM[7714] = MEM[2303] + MEM[3565];
assign MEM[7715] = MEM[2312] + MEM[2313];
assign MEM[7716] = MEM[2324] + MEM[4887];
assign MEM[7717] = MEM[2475] + MEM[3795];
assign MEM[7718] = MEM[2598] + MEM[1039];
assign MEM[7719] = MEM[2643] + MEM[611];
assign MEM[7720] = MEM[2657] + MEM[6422];
assign MEM[7721] = MEM[2671] + MEM[5590];
assign MEM[7722] = MEM[2754] + MEM[342];
assign MEM[7723] = MEM[2844] + MEM[53];
assign MEM[7724] = MEM[2892] + MEM[3330];
assign MEM[7725] = MEM[2899] + MEM[3388];
assign MEM[7726] = MEM[2924] + MEM[3669];
assign MEM[7727] = MEM[2925] + MEM[1445];
assign MEM[7728] = MEM[2974] + MEM[2309];
assign MEM[7729] = MEM[2982] + MEM[826];
assign MEM[7730] = MEM[3012] + MEM[6006];
assign MEM[7731] = MEM[3085] + MEM[4235];
assign MEM[7732] = MEM[3100] + MEM[2287];
assign MEM[7733] = MEM[3122] + MEM[4555];
assign MEM[7734] = MEM[3177] + MEM[3176];
assign MEM[7735] = MEM[3195] + MEM[157];
assign MEM[7736] = MEM[3205] + MEM[4122];
assign MEM[7737] = MEM[3212] + MEM[1941];
assign MEM[7738] = MEM[3228] + MEM[2772];
assign MEM[7739] = MEM[3251] + MEM[5167];
assign MEM[7740] = MEM[3352] + MEM[3353];
assign MEM[7741] = MEM[3354] + MEM[3355];
assign MEM[7742] = MEM[3356] + MEM[7740];
assign MEM[7743] = MEM[3373] + MEM[4364];
assign MEM[7744] = MEM[3441] + MEM[3440];
assign MEM[7745] = MEM[3459] + MEM[5965];
assign MEM[7746] = MEM[3491] + MEM[796];
assign MEM[7747] = MEM[3493] + MEM[5493];
assign MEM[7748] = MEM[3501] + MEM[278];
assign MEM[7749] = MEM[3518] + MEM[2796];
assign MEM[7750] = MEM[3559] + MEM[6196];
assign MEM[7751] = MEM[3592] + MEM[3593];
assign MEM[7752] = MEM[3594] + MEM[3595];
assign MEM[7753] = MEM[3596] + MEM[7751];
assign MEM[7754] = MEM[3628] + MEM[1175];
assign MEM[7755] = MEM[3636] + MEM[574];
assign MEM[7756] = MEM[3667] + MEM[2395];
assign MEM[7757] = MEM[3676] + MEM[4813];
assign MEM[7758] = MEM[3716] + MEM[1506];
assign MEM[7759] = MEM[3779] + MEM[2405];
assign MEM[7760] = MEM[3800] + MEM[3801];
assign MEM[7761] = MEM[3832] + MEM[3833];
assign MEM[7762] = MEM[3839] + MEM[391];
assign MEM[7763] = MEM[3861] + MEM[2315];
assign MEM[7764] = MEM[3875] + MEM[3998];
assign MEM[7765] = MEM[3899] + MEM[6490];
assign MEM[7766] = MEM[3902] + MEM[1374];
assign MEM[7767] = MEM[3979] + MEM[3589];
assign MEM[7768] = MEM[3996] + MEM[3693];
assign MEM[7769] = MEM[4004] + MEM[618];
assign MEM[7770] = MEM[4007] + MEM[6227];
assign MEM[7771] = MEM[4008] + MEM[4009];
assign MEM[7772] = MEM[4015] + MEM[3566];
assign MEM[7773] = MEM[4086] + MEM[750];
assign MEM[7774] = MEM[4143] + MEM[383];
assign MEM[7775] = MEM[4176] + MEM[4177];
assign MEM[7776] = MEM[4264] + MEM[4265];
assign MEM[7777] = MEM[4266] + MEM[4267];
assign MEM[7778] = MEM[4287] + MEM[6155];
assign MEM[7779] = MEM[4346] + MEM[1191];
assign MEM[7780] = MEM[4373] + MEM[4835];
assign MEM[7781] = MEM[4408] + MEM[4409];
assign MEM[7782] = MEM[4418] + MEM[4843];
assign MEM[7783] = MEM[4443] + MEM[3015];
assign MEM[7784] = MEM[4444] + MEM[4515];
assign MEM[7785] = MEM[4451] + MEM[3922];
assign MEM[7786] = MEM[4491] + MEM[5435];
assign MEM[7787] = MEM[4498] + MEM[3428];
assign MEM[7788] = MEM[4512] + MEM[4513];
assign MEM[7789] = MEM[4568] + MEM[4569];
assign MEM[7790] = MEM[4577] + MEM[4576];
assign MEM[7791] = MEM[4585] + MEM[7542];
assign MEM[7792] = MEM[4591] + MEM[421];
assign MEM[7793] = MEM[4593] + MEM[7543];
assign MEM[7794] = MEM[4614] + MEM[4677];
assign MEM[7795] = MEM[4618] + MEM[7319];
assign MEM[7796] = MEM[4647] + MEM[4092];
assign MEM[7797] = MEM[4728] + MEM[4729];
assign MEM[7798] = MEM[4739] + MEM[2750];
assign MEM[7799] = MEM[4799] + MEM[3580];
assign MEM[7800] = MEM[4837] + MEM[1588];
assign MEM[7801] = MEM[4856] + MEM[4857];
assign MEM[7802] = MEM[4871] + MEM[679];
assign MEM[7803] = MEM[4875] + MEM[5643];
assign MEM[7804] = MEM[4904] + MEM[4905];
assign MEM[7805] = MEM[4951] + MEM[4634];
assign MEM[7806] = MEM[4964] + MEM[6330];
assign MEM[7807] = MEM[5032] + MEM[5033];
assign MEM[7808] = MEM[5040] + MEM[5041];
assign MEM[7809] = MEM[5070] + MEM[1711];
assign MEM[7810] = MEM[5090] + MEM[7030];
assign MEM[7811] = MEM[5103] + MEM[2134];
assign MEM[7812] = MEM[5134] + MEM[1494];
assign MEM[7813] = MEM[5183] + MEM[3870];
assign MEM[7814] = MEM[5240] + MEM[5241];
assign MEM[7815] = MEM[5248] + MEM[5249];
assign MEM[7816] = MEM[5256] + MEM[5257];
assign MEM[7817] = MEM[5274] + MEM[7336];
assign MEM[7818] = MEM[5322] + MEM[1622];
assign MEM[7819] = MEM[5330] + MEM[1590];
assign MEM[7820] = MEM[5365] + MEM[47];
assign MEM[7821] = MEM[5384] + MEM[5385];
assign MEM[7822] = MEM[5386] + MEM[5387];
assign MEM[7823] = MEM[5388] + MEM[7821];
assign MEM[7824] = MEM[5402] + MEM[6378];
assign MEM[7825] = MEM[5453] + MEM[842];
assign MEM[7826] = MEM[5468] + MEM[1994];
assign MEM[7827] = MEM[5484] + MEM[31];
assign MEM[7828] = MEM[5491] + MEM[4846];
assign MEM[7829] = MEM[5584] + MEM[5585];
assign MEM[7830] = MEM[5586] + MEM[5587];
assign MEM[7831] = MEM[5588] + MEM[7829];
assign MEM[7832] = MEM[5592] + MEM[5593];
assign MEM[7833] = MEM[5594] + MEM[5595];
assign MEM[7834] = MEM[5596] + MEM[7832];
assign MEM[7835] = MEM[5605] + MEM[3053];
assign MEM[7836] = MEM[5631] + MEM[5789];
assign MEM[7837] = MEM[5636] + MEM[1258];
assign MEM[7838] = MEM[5662] + MEM[5837];
assign MEM[7839] = MEM[5669] + MEM[3187];
assign MEM[7840] = MEM[5677] + MEM[653];
assign MEM[7841] = MEM[5696] + MEM[5697];
assign MEM[7842] = MEM[5704] + MEM[5705];
assign MEM[7843] = MEM[5713] + MEM[5712];
assign MEM[7844] = MEM[5734] + MEM[2756];
assign MEM[7845] = MEM[5749] + MEM[2343];
assign MEM[7846] = MEM[5778] + MEM[5463];
assign MEM[7847] = MEM[5829] + MEM[2039];
assign MEM[7848] = MEM[5846] + MEM[3548];
assign MEM[7849] = MEM[5863] + MEM[839];
assign MEM[7850] = MEM[5915] + MEM[4573];
assign MEM[7851] = MEM[5948] + MEM[4158];
assign MEM[7852] = MEM[5950] + MEM[3277];
assign MEM[7853] = MEM[6008] + MEM[6009];
assign MEM[7854] = MEM[6010] + MEM[7853];
assign MEM[7855] = MEM[6104] + MEM[6105];
assign MEM[7856] = MEM[6106] + MEM[7855];
assign MEM[7857] = MEM[6171] + MEM[4948];
assign MEM[7858] = MEM[6204] + MEM[2659];
assign MEM[7859] = MEM[6207] + MEM[4543];
assign MEM[7860] = MEM[6326] + MEM[6419];
assign MEM[7861] = MEM[6327] + MEM[2279];
assign MEM[7862] = MEM[6329] + MEM[4773];
assign MEM[7863] = MEM[6336] + MEM[6343];
assign MEM[7864] = MEM[6342] + MEM[359];
assign MEM[7865] = MEM[6358] + MEM[584];
assign MEM[7866] = MEM[6360] + MEM[3694];
assign MEM[7867] = MEM[6379] + MEM[6496];
assign MEM[7868] = MEM[6380] + MEM[111];
assign MEM[7869] = MEM[6386] + MEM[6489];
assign MEM[7870] = MEM[6402] + MEM[3453];
assign MEM[7871] = MEM[6440] + MEM[5355];
assign MEM[7872] = MEM[6487] + MEM[93];
assign MEM[7873] = MEM[6499] + MEM[4531];
assign MEM[7874] = MEM[6567] + MEM[2738];
assign MEM[7875] = MEM[7635] + MEM[7636];
assign MEM[7876] = MEM[7638] + MEM[7639];
assign MEM[7877] = MEM[7641] + MEM[7642];
assign MEM[7878] = MEM[7666] + MEM[7667];
assign MEM[7879] = MEM[7682] + MEM[1274];
assign MEM[7880] = MEM[7741] + MEM[7742];
assign MEM[7881] = MEM[7752] + MEM[7753];
assign MEM[7882] = MEM[7776] + MEM[7777];
assign MEM[7883] = MEM[7807] + MEM[5034];
assign MEM[7884] = MEM[7814] + MEM[5242];
assign MEM[7885] = MEM[7815] + MEM[5250];
assign MEM[7886] = MEM[7822] + MEM[7823];
assign MEM[7887] = MEM[7830] + MEM[7831];
assign MEM[7888] = MEM[7833] + MEM[7834];
assign MEM[7889] = MEM[77] + MEM[1315];
assign MEM[7890] = MEM[94] + MEM[3405];
assign MEM[7891] = MEM[173] + MEM[5271];
assign MEM[7892] = MEM[221] + MEM[5196];
assign MEM[7893] = MEM[256] + MEM[257];
assign MEM[7894] = MEM[258] + MEM[259];
assign MEM[7895] = MEM[260] + MEM[7893];
assign MEM[7896] = MEM[320] + MEM[321];
assign MEM[7897] = MEM[326] + MEM[2418];
assign MEM[7898] = MEM[349] + MEM[4172];
assign MEM[7899] = MEM[354] + MEM[1067];
assign MEM[7900] = MEM[358] + MEM[1949];
assign MEM[7901] = MEM[363] + MEM[1298];
assign MEM[7902] = MEM[378] + MEM[5909];
assign MEM[7903] = MEM[389] + MEM[3382];
assign MEM[7904] = MEM[431] + MEM[5349];
assign MEM[7905] = MEM[472] + MEM[473];
assign MEM[7906] = MEM[474] + MEM[475];
assign MEM[7907] = MEM[476] + MEM[7905];
assign MEM[7908] = MEM[578] + MEM[771];
assign MEM[7909] = MEM[579] + MEM[3645];
assign MEM[7910] = MEM[725] + MEM[2871];
assign MEM[7911] = MEM[731] + MEM[843];
assign MEM[7912] = MEM[758] + MEM[4318];
assign MEM[7913] = MEM[760] + MEM[4229];
assign MEM[7914] = MEM[765] + MEM[3886];
assign MEM[7915] = MEM[770] + MEM[2991];
assign MEM[7916] = MEM[820] + MEM[938];
assign MEM[7917] = MEM[821] + MEM[989];
assign MEM[7918] = MEM[822] + MEM[2877];
assign MEM[7919] = MEM[847] + MEM[1228];
assign MEM[7920] = MEM[861] + MEM[1853];
assign MEM[7921] = MEM[928] + MEM[929];
assign MEM[7922] = MEM[949] + MEM[1155];
assign MEM[7923] = MEM[965] + MEM[1077];
assign MEM[7924] = MEM[1024] + MEM[1025];
assign MEM[7925] = MEM[1054] + MEM[1758];
assign MEM[7926] = MEM[1078] + MEM[4500];
assign MEM[7927] = MEM[1096] + MEM[1097];
assign MEM[7928] = MEM[1141] + MEM[4428];
assign MEM[7929] = MEM[1176] + MEM[1177];
assign MEM[7930] = MEM[1236] + MEM[3822];
assign MEM[7931] = MEM[1245] + MEM[38];
assign MEM[7932] = MEM[1295] + MEM[4398];
assign MEM[7933] = MEM[1303] + MEM[3972];
assign MEM[7934] = MEM[1344] + MEM[1345];
assign MEM[7935] = MEM[1346] + MEM[1347];
assign MEM[7936] = MEM[1348] + MEM[7934];
assign MEM[7937] = MEM[1396] + MEM[1986];
assign MEM[7938] = MEM[1434] + MEM[7446];
assign MEM[7939] = MEM[1439] + MEM[2071];
assign MEM[7940] = MEM[1455] + MEM[6203];
assign MEM[7941] = MEM[1466] + MEM[5742];
assign MEM[7942] = MEM[1484] + MEM[1190];
assign MEM[7943] = MEM[1516] + MEM[814];
assign MEM[7944] = MEM[1545] + MEM[1544];
assign MEM[7945] = MEM[1547] + MEM[6376];
assign MEM[7946] = MEM[1599] + MEM[2365];
assign MEM[7947] = MEM[1621] + MEM[5338];
assign MEM[7948] = MEM[1626] + MEM[766];
assign MEM[7949] = MEM[1719] + MEM[3534];
assign MEM[7950] = MEM[1745] + MEM[1744];
assign MEM[7951] = MEM[1762] + MEM[1790];
assign MEM[7952] = MEM[1775] + MEM[3367];
assign MEM[7953] = MEM[1792] + MEM[1793];
assign MEM[7954] = MEM[1794] + MEM[1795];
assign MEM[7955] = MEM[1796] + MEM[7953];
assign MEM[7956] = MEM[1843] + MEM[2661];
assign MEM[7957] = MEM[1958] + MEM[4388];
assign MEM[7958] = MEM[2002] + MEM[5298];
assign MEM[7959] = MEM[2028] + MEM[3821];
assign MEM[7960] = MEM[2058] + MEM[4310];
assign MEM[7961] = MEM[2153] + MEM[2152];
assign MEM[7962] = MEM[2155] + MEM[1877];
assign MEM[7963] = MEM[2169] + MEM[2168];
assign MEM[7964] = MEM[2190] + MEM[143];
assign MEM[7965] = MEM[2224] + MEM[2225];
assign MEM[7966] = MEM[2307] + MEM[2709];
assign MEM[7967] = MEM[2385] + MEM[2384];
assign MEM[7968] = MEM[2413] + MEM[4493];
assign MEM[7969] = MEM[2445] + MEM[4966];
assign MEM[7970] = MEM[2450] + MEM[6426];
assign MEM[7971] = MEM[2463] + MEM[597];
assign MEM[7972] = MEM[2493] + MEM[4525];
assign MEM[7973] = MEM[2535] + MEM[2957];
assign MEM[7974] = MEM[2556] + MEM[1703];
assign MEM[7975] = MEM[2623] + MEM[1419];
assign MEM[7976] = MEM[2653] + MEM[1507];
assign MEM[7977] = MEM[2725] + MEM[5060];
assign MEM[7978] = MEM[2742] + MEM[2622];
assign MEM[7979] = MEM[2778] + MEM[1127];
assign MEM[7980] = MEM[2821] + MEM[5747];
assign MEM[7981] = MEM[2842] + MEM[6505];
assign MEM[7982] = MEM[2859] + MEM[406];
assign MEM[7983] = MEM[2886] + MEM[798];
assign MEM[7984] = MEM[2956] + MEM[3615];
assign MEM[7985] = MEM[2959] + MEM[4452];
assign MEM[7986] = MEM[2998] + MEM[1927];
assign MEM[7987] = MEM[3058] + MEM[3274];
assign MEM[7988] = MEM[3062] + MEM[4095];
assign MEM[7989] = MEM[3091] + MEM[1861];
assign MEM[7990] = MEM[3152] + MEM[3153];
assign MEM[7991] = MEM[3154] + MEM[3155];
assign MEM[7992] = MEM[3182] + MEM[2547];
assign MEM[7993] = MEM[3204] + MEM[3238];
assign MEM[7994] = MEM[3339] + MEM[871];
assign MEM[7995] = MEM[3399] + MEM[3742];
assign MEM[7996] = MEM[3451] + MEM[3450];
assign MEM[7997] = MEM[3487] + MEM[5363];
assign MEM[7998] = MEM[3490] + MEM[6002];
assign MEM[7999] = MEM[3515] + MEM[5114];
assign MEM[8000] = MEM[3573] + MEM[1559];
assign MEM[8001] = MEM[3582] + MEM[3619];
assign MEM[8002] = MEM[3646] + MEM[4807];
assign MEM[8003] = MEM[3715] + MEM[955];
assign MEM[8004] = MEM[3733] + MEM[3789];
assign MEM[8005] = MEM[3751] + MEM[4379];
assign MEM[8006] = MEM[3765] + MEM[1875];
assign MEM[8007] = MEM[3790] + MEM[759];
assign MEM[8008] = MEM[3836] + MEM[3923];
assign MEM[8009] = MEM[3837] + MEM[4348];
assign MEM[8010] = MEM[3853] + MEM[1399];
assign MEM[8011] = MEM[3862] + MEM[5253];
assign MEM[8012] = MEM[3863] + MEM[3571];
assign MEM[8013] = MEM[3895] + MEM[2325];
assign MEM[8014] = MEM[3965] + MEM[1606];
assign MEM[8015] = MEM[3980] + MEM[4596];
assign MEM[8016] = MEM[3997] + MEM[2774];
assign MEM[8017] = MEM[4047] + MEM[3470];
assign MEM[8018] = MEM[4078] + MEM[2694];
assign MEM[8019] = MEM[4082] + MEM[4732];
assign MEM[8020] = MEM[4115] + MEM[1164];
assign MEM[8021] = MEM[4119] + MEM[4579];
assign MEM[8022] = MEM[4136] + MEM[4137];
assign MEM[8023] = MEM[4155] + MEM[5141];
assign MEM[8024] = MEM[4164] + MEM[1493];
assign MEM[8025] = MEM[4173] + MEM[919];
assign MEM[8026] = MEM[4188] + MEM[1062];
assign MEM[8027] = MEM[4199] + MEM[2739];
assign MEM[8028] = MEM[4248] + MEM[4249];
assign MEM[8029] = MEM[4271] + MEM[508];
assign MEM[8030] = MEM[4291] + MEM[3906];
assign MEM[8031] = MEM[4339] + MEM[4652];
assign MEM[8032] = MEM[4499] + MEM[1271];
assign MEM[8033] = MEM[4504] + MEM[4505];
assign MEM[8034] = MEM[4534] + MEM[5884];
assign MEM[8035] = MEM[4536] + MEM[4537];
assign MEM[8036] = MEM[4548] + MEM[1282];
assign MEM[8037] = MEM[4560] + MEM[4561];
assign MEM[8038] = MEM[4606] + MEM[2267];
assign MEM[8039] = MEM[4624] + MEM[4625];
assign MEM[8040] = MEM[4671] + MEM[4684];
assign MEM[8041] = MEM[4701] + MEM[4628];
assign MEM[8042] = MEM[4712] + MEM[4713];
assign MEM[8043] = MEM[4714] + MEM[8042];
assign MEM[8044] = MEM[4766] + MEM[622];
assign MEM[8045] = MEM[4827] + MEM[4826];
assign MEM[8046] = MEM[4851] + MEM[3420];
assign MEM[8047] = MEM[4912] + MEM[4913];
assign MEM[8048] = MEM[4914] + MEM[8047];
assign MEM[8049] = MEM[4960] + MEM[4961];
assign MEM[8050] = MEM[5046] + MEM[3038];
assign MEM[8051] = MEM[5055] + MEM[1014];
assign MEM[8052] = MEM[5066] + MEM[7331];
assign MEM[8053] = MEM[5208] + MEM[5209];
assign MEM[8054] = MEM[5216] + MEM[5217];
assign MEM[8055] = MEM[5232] + MEM[5233];
assign MEM[8056] = MEM[5258] + MEM[7816];
assign MEM[8057] = MEM[5260] + MEM[3011];
assign MEM[8058] = MEM[5302] + MEM[5428];
assign MEM[8059] = MEM[5340] + MEM[3229];
assign MEM[8060] = MEM[5390] + MEM[1090];
assign MEM[8061] = MEM[5391] + MEM[4054];
assign MEM[8062] = MEM[5399] + MEM[125];
assign MEM[8063] = MEM[5411] + MEM[751];
assign MEM[8064] = MEM[5425] + MEM[5424];
assign MEM[8065] = MEM[5431] + MEM[1390];
assign MEM[8066] = MEM[5497] + MEM[5496];
assign MEM[8067] = MEM[5570] + MEM[5975];
assign MEM[8068] = MEM[5575] + MEM[2437];
assign MEM[8069] = MEM[5581] + MEM[1926];
assign MEM[8070] = MEM[5634] + MEM[1357];
assign MEM[8071] = MEM[5679] + MEM[2996];
assign MEM[8072] = MEM[5686] + MEM[463];
assign MEM[8073] = MEM[5716] + MEM[5180];
assign MEM[8074] = MEM[5717] + MEM[2614];
assign MEM[8075] = MEM[5719] + MEM[4390];
assign MEM[8076] = MEM[5725] + MEM[5885];
assign MEM[8077] = MEM[5731] + MEM[2630];
assign MEM[8078] = MEM[5753] + MEM[5752];
assign MEM[8079] = MEM[5780] + MEM[3772];
assign MEM[8080] = MEM[5798] + MEM[1172];
assign MEM[8081] = MEM[5858] + MEM[2851];
assign MEM[8082] = MEM[5867] + MEM[6119];
assign MEM[8083] = MEM[5918] + MEM[638];
assign MEM[8084] = MEM[5952] + MEM[6605];
assign MEM[8085] = MEM[5966] + MEM[3530];
assign MEM[8086] = MEM[6021] + MEM[119];
assign MEM[8087] = MEM[6063] + MEM[1763];
assign MEM[8088] = MEM[6108] + MEM[895];
assign MEM[8089] = MEM[6219] + MEM[962];
assign MEM[8090] = MEM[6247] + MEM[2711];
assign MEM[8091] = MEM[6253] + MEM[5047];
assign MEM[8092] = MEM[6264] + MEM[6265];
assign MEM[8093] = MEM[6266] + MEM[6267];
assign MEM[8094] = MEM[6268] + MEM[8092];
assign MEM[8095] = MEM[6324] + MEM[828];
assign MEM[8096] = MEM[6354] + MEM[1788];
assign MEM[8097] = MEM[6361] + MEM[2263];
assign MEM[8098] = MEM[6365] + MEM[5126];
assign MEM[8099] = MEM[6371] + MEM[903];
assign MEM[8100] = MEM[6385] + MEM[6580];
assign MEM[8101] = MEM[6388] + MEM[6228];
assign MEM[8102] = MEM[6389] + MEM[2452];
assign MEM[8103] = MEM[6390] + MEM[1542];
assign MEM[8104] = MEM[6391] + MEM[2389];
assign MEM[8105] = MEM[6404] + MEM[916];
assign MEM[8106] = MEM[6405] + MEM[836];
assign MEM[8107] = MEM[6409] + MEM[3172];
assign MEM[8108] = MEM[6411] + MEM[6435];
assign MEM[8109] = MEM[6412] + MEM[6414];
assign MEM[8110] = MEM[6418] + MEM[6474];
assign MEM[8111] = MEM[6420] + MEM[6818];
assign MEM[8112] = MEM[6424] + MEM[2403];
assign MEM[8113] = MEM[6429] + MEM[1461];
assign MEM[8114] = MEM[6430] + MEM[4170];
assign MEM[8115] = MEM[6431] + MEM[6500];
assign MEM[8116] = MEM[6433] + MEM[5860];
assign MEM[8117] = MEM[6434] + MEM[5964];
assign MEM[8118] = MEM[6438] + MEM[4946];
assign MEM[8119] = MEM[6442] + MEM[3319];
assign MEM[8120] = MEM[6472] + MEM[5628];
assign MEM[8121] = MEM[6477] + MEM[2492];
assign MEM[8122] = MEM[6478] + MEM[6004];
assign MEM[8123] = MEM[6491] + MEM[3579];
assign MEM[8124] = MEM[6497] + MEM[4203];
assign MEM[8125] = MEM[6501] + MEM[3918];
assign MEM[8126] = MEM[6506] + MEM[6507];
assign MEM[8127] = MEM[6581] + MEM[3658];
assign MEM[8128] = MEM[6592] + MEM[6436];
assign MEM[8129] = MEM[6634] + MEM[6464];
assign MEM[8130] = MEM[6636] + MEM[738];
assign MEM[8131] = MEM[6650] + MEM[6651];
assign MEM[8132] = MEM[6722] + MEM[6598];
assign MEM[8133] = MEM[6742] + MEM[6538];
assign MEM[8134] = MEM[6855] + MEM[1810];
assign MEM[8135] = MEM[6947] + MEM[1314];
assign MEM[8136] = MEM[7333] + MEM[5226];
assign MEM[8137] = MEM[7894] + MEM[7895];
assign MEM[8138] = MEM[7896] + MEM[322];
assign MEM[8139] = MEM[7906] + MEM[7907];
assign MEM[8140] = MEM[7921] + MEM[930];
assign MEM[8141] = MEM[7935] + MEM[7936];
assign MEM[8142] = MEM[7954] + MEM[7955];
assign MEM[8143] = MEM[7990] + MEM[7991];
assign MEM[8144] = MEM[7996] + MEM[6577];
assign MEM[8145] = MEM[8039] + MEM[4626];
assign MEM[8146] = MEM[8093] + MEM[8094];
assign MEM[8147] = MEM[8114] + MEM[6587];
assign MEM[8148] = MEM[30] + MEM[1154];
assign MEM[8149] = MEM[101] + MEM[886];
assign MEM[8150] = MEM[112] + MEM[113];
assign MEM[8151] = MEM[114] + MEM[115];
assign MEM[8152] = MEM[128] + MEM[129];
assign MEM[8153] = MEM[130] + MEM[131];
assign MEM[8154] = MEM[132] + MEM[8152];
assign MEM[8155] = MEM[165] + MEM[246];
assign MEM[8156] = MEM[176] + MEM[177];
assign MEM[8157] = MEM[178] + MEM[179];
assign MEM[8158] = MEM[180] + MEM[8156];
assign MEM[8159] = MEM[207] + MEM[1671];
assign MEM[8160] = MEM[237] + MEM[2116];
assign MEM[8161] = MEM[238] + MEM[5404];
assign MEM[8162] = MEM[286] + MEM[413];
assign MEM[8163] = MEM[307] + MEM[3219];
assign MEM[8164] = MEM[331] + MEM[478];
assign MEM[8165] = MEM[334] + MEM[373];
assign MEM[8166] = MEM[338] + MEM[1731];
assign MEM[8167] = MEM[339] + MEM[3686];
assign MEM[8168] = MEM[366] + MEM[1242];
assign MEM[8169] = MEM[372] + MEM[3157];
assign MEM[8170] = MEM[390] + MEM[471];
assign MEM[8171] = MEM[411] + MEM[1594];
assign MEM[8172] = MEM[415] + MEM[2283];
assign MEM[8173] = MEM[430] + MEM[715];
assign MEM[8174] = MEM[477] + MEM[2123];
assign MEM[8175] = MEM[500] + MEM[3934];
assign MEM[8176] = MEM[549] + MEM[3446];
assign MEM[8177] = MEM[554] + MEM[1444];
assign MEM[8178] = MEM[563] + MEM[1156];
assign MEM[8179] = MEM[564] + MEM[3115];
assign MEM[8180] = MEM[604] + MEM[4011];
assign MEM[8181] = MEM[621] + MEM[5814];
assign MEM[8182] = MEM[678] + MEM[943];
assign MEM[8183] = MEM[685] + MEM[2340];
assign MEM[8184] = MEM[732] + MEM[3735];
assign MEM[8185] = MEM[733] + MEM[730];
assign MEM[8186] = MEM[762] + MEM[6029];
assign MEM[8187] = MEM[763] + MEM[2890];
assign MEM[8188] = MEM[772] + MEM[95];
assign MEM[8189] = MEM[774] + MEM[2029];
assign MEM[8190] = MEM[777] + MEM[776];
assign MEM[8191] = MEM[785] + MEM[784];
assign MEM[8192] = MEM[804] + MEM[2142];
assign MEM[8193] = MEM[807] + MEM[4403];
assign MEM[8194] = MEM[859] + MEM[2775];
assign MEM[8195] = MEM[879] + MEM[1358];
assign MEM[8196] = MEM[904] + MEM[905];
assign MEM[8197] = MEM[906] + MEM[907];
assign MEM[8198] = MEM[908] + MEM[8196];
assign MEM[8199] = MEM[934] + MEM[3852];
assign MEM[8200] = MEM[948] + MEM[1082];
assign MEM[8201] = MEM[964] + MEM[1915];
assign MEM[8202] = MEM[971] + MEM[4075];
assign MEM[8203] = MEM[984] + MEM[985];
assign MEM[8204] = MEM[997] + MEM[571];
assign MEM[8205] = MEM[1001] + MEM[1000];
assign MEM[8206] = MEM[1021] + MEM[1142];
assign MEM[8207] = MEM[1028] + MEM[3331];
assign MEM[8208] = MEM[1066] + MEM[5462];
assign MEM[8209] = MEM[1079] + MEM[2382];
assign MEM[8210] = MEM[1143] + MEM[935];
assign MEM[8211] = MEM[1223] + MEM[2135];
assign MEM[8212] = MEM[1226] + MEM[7085];
assign MEM[8213] = MEM[1238] + MEM[2855];
assign MEM[8214] = MEM[1250] + MEM[7680];
assign MEM[8215] = MEM[1267] + MEM[6214];
assign MEM[8216] = MEM[1349] + MEM[6199];
assign MEM[8217] = MEM[1422] + MEM[4762];
assign MEM[8218] = MEM[1426] + MEM[3412];
assign MEM[8219] = MEM[1467] + MEM[2710];
assign MEM[8220] = MEM[1490] + MEM[3315];
assign MEM[8221] = MEM[1549] + MEM[5091];
assign MEM[8222] = MEM[1551] + MEM[4658];
assign MEM[8223] = MEM[1563] + MEM[1670];
assign MEM[8224] = MEM[1576] + MEM[1577];
assign MEM[8225] = MEM[1647] + MEM[3222];
assign MEM[8226] = MEM[1656] + MEM[1657];
assign MEM[8227] = MEM[1683] + MEM[6115];
assign MEM[8228] = MEM[1734] + MEM[2252];
assign MEM[8229] = MEM[1818] + MEM[5159];
assign MEM[8230] = MEM[1826] + MEM[4062];
assign MEM[8231] = MEM[1827] + MEM[4334];
assign MEM[8232] = MEM[1844] + MEM[1495];
assign MEM[8233] = MEM[1876] + MEM[2333];
assign MEM[8234] = MEM[1878] + MEM[3046];
assign MEM[8235] = MEM[1932] + MEM[3044];
assign MEM[8236] = MEM[1936] + MEM[1937];
assign MEM[8237] = MEM[1959] + MEM[5939];
assign MEM[8238] = MEM[1991] + MEM[1477];
assign MEM[8239] = MEM[2046] + MEM[3590];
assign MEM[8240] = MEM[2069] + MEM[4354];
assign MEM[8241] = MEM[2083] + MEM[3604];
assign MEM[8242] = MEM[2124] + MEM[1510];
assign MEM[8243] = MEM[2148] + MEM[1838];
assign MEM[8244] = MEM[2150] + MEM[3478];
assign MEM[8245] = MEM[2188] + MEM[4750];
assign MEM[8246] = MEM[2223] + MEM[1045];
assign MEM[8247] = MEM[2247] + MEM[3350];
assign MEM[8248] = MEM[2284] + MEM[3591];
assign MEM[8249] = MEM[2332] + MEM[2342];
assign MEM[8250] = MEM[2347] + MEM[4220];
assign MEM[8251] = MEM[2371] + MEM[4430];
assign MEM[8252] = MEM[2383] + MEM[3829];
assign MEM[8253] = MEM[2411] + MEM[1651];
assign MEM[8254] = MEM[2435] + MEM[1269];
assign MEM[8255] = MEM[2439] + MEM[1284];
assign MEM[8256] = MEM[2460] + MEM[1940];
assign MEM[8257] = MEM[2499] + MEM[3527];
assign MEM[8258] = MEM[2509] + MEM[3956];
assign MEM[8259] = MEM[2516] + MEM[1831];
assign MEM[8260] = MEM[2526] + MEM[261];
assign MEM[8261] = MEM[2539] + MEM[4276];
assign MEM[8262] = MEM[2543] + MEM[4391];
assign MEM[8263] = MEM[2582] + MEM[1402];
assign MEM[8264] = MEM[2762] + MEM[2782];
assign MEM[8265] = MEM[2829] + MEM[1100];
assign MEM[8266] = MEM[2836] + MEM[1885];
assign MEM[8267] = MEM[2858] + MEM[2118];
assign MEM[8268] = MEM[2885] + MEM[2189];
assign MEM[8269] = MEM[2898] + MEM[1556];
assign MEM[8270] = MEM[2910] + MEM[2053];
assign MEM[8271] = MEM[3022] + MEM[1582];
assign MEM[8272] = MEM[3076] + MEM[6415];
assign MEM[8273] = MEM[3099] + MEM[2780];
assign MEM[8274] = MEM[3117] + MEM[4810];
assign MEM[8275] = MEM[3123] + MEM[4866];
assign MEM[8276] = MEM[3133] + MEM[5622];
assign MEM[8277] = MEM[3151] + MEM[802];
assign MEM[8278] = MEM[3253] + MEM[3917];
assign MEM[8279] = MEM[3263] + MEM[5434];
assign MEM[8280] = MEM[3264] + MEM[3265];
assign MEM[8281] = MEM[3403] + MEM[6578];
assign MEM[8282] = MEM[3436] + MEM[332];
assign MEM[8283] = MEM[3460] + MEM[6480];
assign MEM[8284] = MEM[3466] + MEM[3474];
assign MEM[8285] = MEM[3475] + MEM[4221];
assign MEM[8286] = MEM[3522] + MEM[5044];
assign MEM[8287] = MEM[3524] + MEM[6463];
assign MEM[8288] = MEM[3554] + MEM[2986];
assign MEM[8289] = MEM[3564] + MEM[4251];
assign MEM[8290] = MEM[3652] + MEM[6116];
assign MEM[8291] = MEM[3653] + MEM[5429];
assign MEM[8292] = MEM[3675] + MEM[3627];
assign MEM[8293] = MEM[3701] + MEM[4803];
assign MEM[8294] = MEM[3709] + MEM[429];
assign MEM[8295] = MEM[3717] + MEM[3181];
assign MEM[8296] = MEM[3731] + MEM[2963];
assign MEM[8297] = MEM[3774] + MEM[3413];
assign MEM[8298] = MEM[3778] + MEM[4130];
assign MEM[8299] = MEM[3842] + MEM[1085];
assign MEM[8300] = MEM[3946] + MEM[3754];
assign MEM[8301] = MEM[3994] + MEM[4419];
assign MEM[8302] = MEM[4094] + MEM[893];
assign MEM[8303] = MEM[4108] + MEM[3477];
assign MEM[8304] = MEM[4140] + MEM[1685];
assign MEM[8305] = MEM[4247] + MEM[894];
assign MEM[8306] = MEM[4288] + MEM[4289];
assign MEM[8307] = MEM[4333] + MEM[2215];
assign MEM[8308] = MEM[4471] + MEM[2951];
assign MEM[8309] = MEM[4502] + MEM[2530];
assign MEM[8310] = MEM[4582] + MEM[4526];
assign MEM[8311] = MEM[4588] + MEM[5455];
assign MEM[8312] = MEM[4595] + MEM[4421];
assign MEM[8313] = MEM[4605] + MEM[5358];
assign MEM[8314] = MEM[4620] + MEM[340];
assign MEM[8315] = MEM[4630] + MEM[6023];
assign MEM[8316] = MEM[4636] + MEM[5158];
assign MEM[8317] = MEM[4670] + MEM[4818];
assign MEM[8318] = MEM[4759] + MEM[5245];
assign MEM[8319] = MEM[4795] + MEM[2447];
assign MEM[8320] = MEM[4804] + MEM[3551];
assign MEM[8321] = MEM[4874] + MEM[4639];
assign MEM[8322] = MEM[4918] + MEM[5527];
assign MEM[8323] = MEM[4933] + MEM[2021];
assign MEM[8324] = MEM[4973] + MEM[2076];
assign MEM[8325] = MEM[4980] + MEM[783];
assign MEM[8326] = MEM[5068] + MEM[3567];
assign MEM[8327] = MEM[5076] + MEM[5621];
assign MEM[8328] = MEM[5136] + MEM[5137];
assign MEM[8329] = MEM[5138] + MEM[8328];
assign MEM[8330] = MEM[5197] + MEM[2258];
assign MEM[8331] = MEM[5206] + MEM[5052];
assign MEM[8332] = MEM[5237] + MEM[3620];
assign MEM[8333] = MEM[5247] + MEM[2478];
assign MEM[8334] = MEM[5259] + MEM[2908];
assign MEM[8335] = MEM[5277] + MEM[5941];
assign MEM[8336] = MEM[5284] + MEM[55];
assign MEM[8337] = MEM[5292] + MEM[5859];
assign MEM[8338] = MEM[5307] + MEM[5525];
assign MEM[8339] = MEM[5310] + MEM[761];
assign MEM[8340] = MEM[5334] + MEM[634];
assign MEM[8341] = MEM[5368] + MEM[5369];
assign MEM[8342] = MEM[5370] + MEM[5371];
assign MEM[8343] = MEM[5372] + MEM[8341];
assign MEM[8344] = MEM[5382] + MEM[3644];
assign MEM[8345] = MEM[5392] + MEM[5393];
assign MEM[8346] = MEM[5394] + MEM[8345];
assign MEM[8347] = MEM[5427] + MEM[1525];
assign MEM[8348] = MEM[5439] + MEM[4564];
assign MEM[8349] = MEM[5470] + MEM[3626];
assign MEM[8350] = MEM[5472] + MEM[5473];
assign MEM[8351] = MEM[5477] + MEM[1246];
assign MEM[8352] = MEM[5530] + MEM[5275];
assign MEM[8353] = MEM[5540] + MEM[2062];
assign MEM[8354] = MEM[5549] + MEM[2874];
assign MEM[8355] = MEM[5559] + MEM[6471];
assign MEM[8356] = MEM[5646] + MEM[2092];
assign MEM[8357] = MEM[5655] + MEM[662];
assign MEM[8358] = MEM[5668] + MEM[5874];
assign MEM[8359] = MEM[5680] + MEM[5681];
assign MEM[8360] = MEM[5687] + MEM[2197];
assign MEM[8361] = MEM[5743] + MEM[1922];
assign MEM[8362] = MEM[5762] + MEM[2156];
assign MEM[8363] = MEM[5764] + MEM[3931];
assign MEM[8364] = MEM[5787] + MEM[6441];
assign MEM[8365] = MEM[5894] + MEM[2973];
assign MEM[8366] = MEM[5898] + MEM[4085];
assign MEM[8367] = MEM[5931] + MEM[5763];
assign MEM[8368] = MEM[5934] + MEM[2454];
assign MEM[8369] = MEM[5938] + MEM[2114];
assign MEM[8370] = MEM[5943] + MEM[5999];
assign MEM[8371] = MEM[5949] + MEM[1575];
assign MEM[8372] = MEM[5953] + MEM[5954];
assign MEM[8373] = MEM[6072] + MEM[6073];
assign MEM[8374] = MEM[6074] + MEM[6075];
assign MEM[8375] = MEM[6076] + MEM[8373];
assign MEM[8376] = MEM[6139] + MEM[6162];
assign MEM[8377] = MEM[6154] + MEM[2828];
assign MEM[8378] = MEM[6156] + MEM[619];
assign MEM[8379] = MEM[6212] + MEM[3908];
assign MEM[8380] = MEM[6220] + MEM[2749];
assign MEM[8381] = MEM[6416] + MEM[5514];
assign MEM[8382] = MEM[6421] + MEM[2519];
assign MEM[8383] = MEM[6423] + MEM[3098];
assign MEM[8384] = MEM[6427] + MEM[3955];
assign MEM[8385] = MEM[6443] + MEM[3226];
assign MEM[8386] = MEM[6476] + MEM[6546];
assign MEM[8387] = MEM[6485] + MEM[2604];
assign MEM[8388] = MEM[6492] + MEM[4527];
assign MEM[8389] = MEM[6495] + MEM[5507];
assign MEM[8390] = MEM[6512] + MEM[2490];
assign MEM[8391] = MEM[6516] + MEM[5059];
assign MEM[8392] = MEM[6548] + MEM[5082];
assign MEM[8393] = MEM[6557] + MEM[7017];
assign MEM[8394] = MEM[6562] + MEM[3359];
assign MEM[8395] = MEM[6571] + MEM[6575];
assign MEM[8396] = MEM[6576] + MEM[2551];
assign MEM[8397] = MEM[6588] + MEM[374];
assign MEM[8398] = MEM[6606] + MEM[5564];
assign MEM[8399] = MEM[6612] + MEM[507];
assign MEM[8400] = MEM[6637] + MEM[858];
assign MEM[8401] = MEM[6663] + MEM[2130];
assign MEM[8402] = MEM[6673] + MEM[6671];
assign MEM[8403] = MEM[6724] + MEM[6723];
assign MEM[8404] = MEM[6778] + MEM[6784];
assign MEM[8405] = MEM[6802] + MEM[1386];
assign MEM[8406] = MEM[6820] + MEM[2410];
assign MEM[8407] = MEM[8150] + MEM[8151];
assign MEM[8408] = MEM[8153] + MEM[8154];
assign MEM[8409] = MEM[8157] + MEM[8158];
assign MEM[8410] = MEM[8197] + MEM[8198];
assign MEM[8411] = MEM[8342] + MEM[8343];
assign MEM[8412] = MEM[8350] + MEM[5474];
assign MEM[8413] = MEM[8374] + MEM[8375];
assign MEM[8414] = MEM[62] + MEM[4159];
assign MEM[8415] = MEM[86] + MEM[2693];
assign MEM[8416] = MEM[167] + MEM[3683];
assign MEM[8417] = MEM[214] + MEM[2868];
assign MEM[8418] = MEM[230] + MEM[1253];
assign MEM[8419] = MEM[255] + MEM[4039];
assign MEM[8420] = MEM[302] + MEM[2893];
assign MEM[8421] = MEM[464] + MEM[465];
assign MEM[8422] = MEM[466] + MEM[467];
assign MEM[8423] = MEM[468] + MEM[8421];
assign MEM[8424] = MEM[484] + MEM[1412];
assign MEM[8425] = MEM[486] + MEM[3021];
assign MEM[8426] = MEM[519] + MEM[4037];
assign MEM[8427] = MEM[524] + MEM[2301];
assign MEM[8428] = MEM[551] + MEM[1479];
assign MEM[8429] = MEM[575] + MEM[1981];
assign MEM[8430] = MEM[670] + MEM[6662];
assign MEM[8431] = MEM[687] + MEM[1738];
assign MEM[8432] = MEM[718] + MEM[2966];
assign MEM[8433] = MEM[815] + MEM[3170];
assign MEM[8434] = MEM[823] + MEM[2559];
assign MEM[8435] = MEM[850] + MEM[166];
assign MEM[8436] = MEM[876] + MEM[644];
assign MEM[8437] = MEM[915] + MEM[1483];
assign MEM[8438] = MEM[933] + MEM[1487];
assign MEM[8439] = MEM[939] + MEM[2980];
assign MEM[8440] = MEM[976] + MEM[977];
assign MEM[8441] = MEM[1030] + MEM[1371];
assign MEM[8442] = MEM[1060] + MEM[3685];
assign MEM[8443] = MEM[1068] + MEM[3202];
assign MEM[8444] = MEM[1087] + MEM[4431];
assign MEM[8445] = MEM[1093] + MEM[2487];
assign MEM[8446] = MEM[1107] + MEM[2007];
assign MEM[8447] = MEM[1117] + MEM[4327];
assign MEM[8448] = MEM[1135] + MEM[1239];
assign MEM[8449] = MEM[1144] + MEM[1145];
assign MEM[8450] = MEM[1147] + MEM[3051];
assign MEM[8451] = MEM[1167] + MEM[1859];
assign MEM[8452] = MEM[1230] + MEM[3966];
assign MEM[8453] = MEM[1360] + MEM[1361];
assign MEM[8454] = MEM[1362] + MEM[8453];
assign MEM[8455] = MEM[1364] + MEM[3271];
assign MEM[8456] = MEM[1380] + MEM[972];
assign MEM[8457] = MEM[1389] + MEM[6545];
assign MEM[8458] = MEM[1394] + MEM[5045];
assign MEM[8459] = MEM[1403] + MEM[1331];
assign MEM[8460] = MEM[1414] + MEM[3019];
assign MEM[8461] = MEM[1415] + MEM[4343];
assign MEM[8462] = MEM[1428] + MEM[3165];
assign MEM[8463] = MEM[1458] + MEM[1459];
assign MEM[8464] = MEM[1475] + MEM[2391];
assign MEM[8465] = MEM[1514] + MEM[1515];
assign MEM[8466] = MEM[1531] + MEM[5110];
assign MEM[8467] = MEM[1533] + MEM[6879];
assign MEM[8468] = MEM[1558] + MEM[3167];
assign MEM[8469] = MEM[1564] + MEM[2799];
assign MEM[8470] = MEM[1573] + MEM[5508];
assign MEM[8471] = MEM[1620] + MEM[5317];
assign MEM[8472] = MEM[1637] + MEM[5436];
assign MEM[8473] = MEM[1666] + MEM[7696];
assign MEM[8474] = MEM[1667] + MEM[1227];
assign MEM[8475] = MEM[1699] + MEM[2570];
assign MEM[8476] = MEM[1701] + MEM[2285];
assign MEM[8477] = MEM[1740] + MEM[1722];
assign MEM[8478] = MEM[1759] + MEM[2610];
assign MEM[8479] = MEM[1807] + MEM[2388];
assign MEM[8480] = MEM[1850] + MEM[7459];
assign MEM[8481] = MEM[1868] + MEM[3103];
assign MEM[8482] = MEM[1874] + MEM[3398];
assign MEM[8483] = MEM[1890] + MEM[1891];
assign MEM[8484] = MEM[1909] + MEM[3642];
assign MEM[8485] = MEM[1911] + MEM[4023];
assign MEM[8486] = MEM[1923] + MEM[5879];
assign MEM[8487] = MEM[1933] + MEM[5243];
assign MEM[8488] = MEM[1948] + MEM[4509];
assign MEM[8489] = MEM[1975] + MEM[4645];
assign MEM[8490] = MEM[1990] + MEM[5031];
assign MEM[8491] = MEM[2022] + MEM[2571];
assign MEM[8492] = MEM[2043] + MEM[5021];
assign MEM[8493] = MEM[2088] + MEM[2089];
assign MEM[8494] = MEM[2108] + MEM[3611];
assign MEM[8495] = MEM[2119] + MEM[439];
assign MEM[8496] = MEM[2161] + MEM[2160];
assign MEM[8497] = MEM[2204] + MEM[3214];
assign MEM[8498] = MEM[2210] + MEM[4079];
assign MEM[8499] = MEM[2229] + MEM[2228];
assign MEM[8500] = MEM[2236] + MEM[3124];
assign MEM[8501] = MEM[2293] + MEM[2786];
assign MEM[8502] = MEM[2334] + MEM[4293];
assign MEM[8503] = MEM[2349] + MEM[5979];
assign MEM[8504] = MEM[2355] + MEM[4070];
assign MEM[8505] = MEM[2397] + MEM[4211];
assign MEM[8506] = MEM[2446] + MEM[387];
assign MEM[8507] = MEM[2464] + MEM[2465];
assign MEM[8508] = MEM[2466] + MEM[2467];
assign MEM[8509] = MEM[2479] + MEM[3699];
assign MEM[8510] = MEM[2502] + MEM[3276];
assign MEM[8511] = MEM[2525] + MEM[6269];
assign MEM[8512] = MEM[2533] + MEM[2507];
assign MEM[8513] = MEM[2555] + MEM[3983];
assign MEM[8514] = MEM[2597] + MEM[2909];
assign MEM[8515] = MEM[2652] + MEM[2557];
assign MEM[8516] = MEM[2759] + MEM[3071];
assign MEM[8517] = MEM[2831] + MEM[4716];
assign MEM[8518] = MEM[2867] + MEM[4530];
assign MEM[8519] = MEM[2975] + MEM[5124];
assign MEM[8520] = MEM[2990] + MEM[6147];
assign MEM[8521] = MEM[3003] + MEM[3538];
assign MEM[8522] = MEM[3026] + MEM[7284];
assign MEM[8523] = MEM[3060] + MEM[3623];
assign MEM[8524] = MEM[3110] + MEM[3131];
assign MEM[8525] = MEM[3116] + MEM[4003];
assign MEM[8526] = MEM[3125] + MEM[3445];
assign MEM[8527] = MEM[3134] + MEM[126];
assign MEM[8528] = MEM[3162] + MEM[4317];
assign MEM[8529] = MEM[3232] + MEM[3233];
assign MEM[8530] = MEM[3317] + MEM[3989];
assign MEM[8531] = MEM[3379] + MEM[3575];
assign MEM[8532] = MEM[3443] + MEM[3691];
assign MEM[8533] = MEM[3508] + MEM[3942];
assign MEM[8534] = MEM[3542] + MEM[2718];
assign MEM[8535] = MEM[3550] + MEM[6444];
assign MEM[8536] = MEM[3603] + MEM[4150];
assign MEM[8537] = MEM[3622] + MEM[356];
assign MEM[8538] = MEM[3638] + MEM[4805];
assign MEM[8539] = MEM[3708] + MEM[71];
assign MEM[8540] = MEM[3727] + MEM[5533];
assign MEM[8541] = MEM[3740] + MEM[4335];
assign MEM[8542] = MEM[3755] + MEM[5107];
assign MEM[8543] = MEM[3756] + MEM[5755];
assign MEM[8544] = MEM[3782] + MEM[4959];
assign MEM[8545] = MEM[3804] + MEM[4165];
assign MEM[8546] = MEM[3814] + MEM[3334];
assign MEM[8547] = MEM[3827] + MEM[3826];
assign MEM[8548] = MEM[3843] + MEM[4663];
assign MEM[8549] = MEM[3846] + MEM[4994];
assign MEM[8550] = MEM[3884] + MEM[4661];
assign MEM[8551] = MEM[3894] + MEM[3758];
assign MEM[8552] = MEM[3914] + MEM[2061];
assign MEM[8553] = MEM[4030] + MEM[6470];
assign MEM[8554] = MEM[4051] + MEM[6534];
assign MEM[8555] = MEM[4099] + MEM[1935];
assign MEM[8556] = MEM[4239] + MEM[1263];
assign MEM[8557] = MEM[4245] + MEM[5438];
assign MEM[8558] = MEM[4250] + MEM[1266];
assign MEM[8559] = MEM[4269] + MEM[3796];
assign MEM[8560] = MEM[4308] + MEM[3878];
assign MEM[8561] = MEM[4314] + MEM[4315];
assign MEM[8562] = MEM[4319] + MEM[5101];
assign MEM[8563] = MEM[4330] + MEM[4338];
assign MEM[8564] = MEM[4332] + MEM[4863];
assign MEM[8565] = MEM[4355] + MEM[5452];
assign MEM[8566] = MEM[4363] + MEM[5733];
assign MEM[8567] = MEM[4366] + MEM[2727];
assign MEM[8568] = MEM[4399] + MEM[4646];
assign MEM[8569] = MEM[4436] + MEM[3971];
assign MEM[8570] = MEM[4487] + MEM[2277];
assign MEM[8571] = MEM[4518] + MEM[4838];
assign MEM[8572] = MEM[4598] + MEM[717];
assign MEM[8573] = MEM[4612] + MEM[6465];
assign MEM[8574] = MEM[4615] + MEM[4870];
assign MEM[8575] = MEM[4655] + MEM[4738];
assign MEM[8576] = MEM[4662] + MEM[967];
assign MEM[8577] = MEM[4678] + MEM[6523];
assign MEM[8578] = MEM[4735] + MEM[2367];
assign MEM[8579] = MEM[4743] + MEM[5140];
assign MEM[8580] = MEM[4774] + MEM[2415];
assign MEM[8581] = MEM[4778] + MEM[645];
assign MEM[8582] = MEM[4791] + MEM[5460];
assign MEM[8583] = MEM[4820] + MEM[954];
assign MEM[8584] = MEM[4853] + MEM[5142];
assign MEM[8585] = MEM[4908] + MEM[5188];
assign MEM[8586] = MEM[4916] + MEM[4915];
assign MEM[8587] = MEM[4987] + MEM[5724];
assign MEM[8588] = MEM[5020] + MEM[6481];
assign MEM[8589] = MEM[5078] + MEM[3135];
assign MEM[8590] = MEM[5083] + MEM[5524];
assign MEM[8591] = MEM[5149] + MEM[6245];
assign MEM[8592] = MEM[5160] + MEM[5161];
assign MEM[8593] = MEM[5162] + MEM[5163];
assign MEM[8594] = MEM[5164] + MEM[8592];
assign MEM[8595] = MEM[5195] + MEM[5996];
assign MEM[8596] = MEM[5228] + MEM[3871];
assign MEM[8597] = MEM[5231] + MEM[855];
assign MEM[8598] = MEM[5251] + MEM[5951];
assign MEM[8599] = MEM[5269] + MEM[5487];
assign MEM[8600] = MEM[5359] + MEM[4885];
assign MEM[8601] = MEM[5366] + MEM[6563];
assign MEM[8602] = MEM[5373] + MEM[4396];
assign MEM[8603] = MEM[5398] + MEM[6211];
assign MEM[8604] = MEM[5421] + MEM[941];
assign MEM[8605] = MEM[5526] + MEM[740];
assign MEM[8606] = MEM[5538] + MEM[846];
assign MEM[8607] = MEM[5652] + MEM[343];
assign MEM[8608] = MEM[5674] + MEM[6094];
assign MEM[8609] = MEM[5676] + MEM[3973];
assign MEM[8610] = MEM[5691] + MEM[1980];
assign MEM[8611] = MEM[5718] + MEM[1003];
assign MEM[8612] = MEM[5726] + MEM[5318];
assign MEM[8613] = MEM[5727] + MEM[1836];
assign MEM[8614] = MEM[5765] + MEM[2356];
assign MEM[8615] = MEM[5767] + MEM[197];
assign MEM[8616] = MEM[5783] + MEM[5788];
assign MEM[8617] = MEM[5870] + MEM[3077];
assign MEM[8618] = MEM[5887] + MEM[3805];
assign MEM[8619] = MEM[5936] + MEM[2322];
assign MEM[8620] = MEM[5956] + MEM[587];
assign MEM[8621] = MEM[6013] + MEM[447];
assign MEM[8622] = MEM[6038] + MEM[3511];
assign MEM[8623] = MEM[6048] + MEM[6049];
assign MEM[8624] = MEM[6050] + MEM[6051];
assign MEM[8625] = MEM[6052] + MEM[8623];
assign MEM[8626] = MEM[6055] + MEM[2947];
assign MEM[8627] = MEM[6096] + MEM[6097];
assign MEM[8628] = MEM[6098] + MEM[6099];
assign MEM[8629] = MEM[6100] + MEM[8627];
assign MEM[8630] = MEM[6103] + MEM[1610];
assign MEM[8631] = MEM[6125] + MEM[4127];
assign MEM[8632] = MEM[6150] + MEM[6222];
assign MEM[8633] = MEM[6240] + MEM[6241];
assign MEM[8634] = MEM[6242] + MEM[6243];
assign MEM[8635] = MEM[6244] + MEM[8633];
assign MEM[8636] = MEM[6445] + MEM[2213];
assign MEM[8637] = MEM[6446] + MEM[1133];
assign MEM[8638] = MEM[6455] + MEM[6667];
assign MEM[8639] = MEM[6462] + MEM[1429];
assign MEM[8640] = MEM[6468] + MEM[1523];
assign MEM[8641] = MEM[6473] + MEM[2962];
assign MEM[8642] = MEM[6484] + MEM[3700];
assign MEM[8643] = MEM[6486] + MEM[4375];
assign MEM[8644] = MEM[6493] + MEM[6494];
assign MEM[8645] = MEM[6498] + MEM[1925];
assign MEM[8646] = MEM[6513] + MEM[3215];
assign MEM[8647] = MEM[6514] + MEM[1454];
assign MEM[8648] = MEM[6515] + MEM[6175];
assign MEM[8649] = MEM[6517] + MEM[4909];
assign MEM[8650] = MEM[6524] + MEM[6031];
assign MEM[8651] = MEM[6525] + MEM[764];
assign MEM[8652] = MEM[6536] + MEM[546];
assign MEM[8653] = MEM[6555] + MEM[231];
assign MEM[8654] = MEM[6564] + MEM[6716];
assign MEM[8655] = MEM[6565] + MEM[2532];
assign MEM[8656] = MEM[6566] + MEM[3941];
assign MEM[8657] = MEM[6570] + MEM[1335];
assign MEM[8658] = MEM[6583] + MEM[6695];
assign MEM[8659] = MEM[6585] + MEM[15];
assign MEM[8660] = MEM[6589] + MEM[2965];
assign MEM[8661] = MEM[6590] + MEM[3190];
assign MEM[8662] = MEM[6591] + MEM[3900];
assign MEM[8663] = MEM[6593] + MEM[2077];
assign MEM[8664] = MEM[6608] + MEM[6672];
assign MEM[8665] = MEM[6618] + MEM[206];
assign MEM[8666] = MEM[6631] + MEM[6537];
assign MEM[8667] = MEM[6657] + MEM[6963];
assign MEM[8668] = MEM[6668] + MEM[2146];
assign MEM[8669] = MEM[6669] + MEM[2442];
assign MEM[8670] = MEM[6683] + MEM[7128];
assign MEM[8671] = MEM[6686] + MEM[2667];
assign MEM[8672] = MEM[6696] + MEM[1715];
assign MEM[8673] = MEM[6702] + MEM[6854];
assign MEM[8674] = MEM[6708] + MEM[4819];
assign MEM[8675] = MEM[6737] + MEM[4087];
assign MEM[8676] = MEM[6750] + MEM[4437];
assign MEM[8677] = MEM[6798] + MEM[6941];
assign MEM[8678] = MEM[6844] + MEM[6584];
assign MEM[8679] = MEM[6896] + MEM[6699];
assign MEM[8680] = MEM[6956] + MEM[1714];
assign MEM[8681] = MEM[6977] + MEM[6815];
assign MEM[8682] = MEM[6994] + MEM[6582];
assign MEM[8683] = MEM[7033] + MEM[5410];
assign MEM[8684] = MEM[8422] + MEM[8423];
assign MEM[8685] = MEM[8449] + MEM[1146];
assign MEM[8686] = MEM[8483] + MEM[6960];
assign MEM[8687] = MEM[8507] + MEM[8508];
assign MEM[8688] = MEM[8547] + MEM[7303];
assign MEM[8689] = MEM[8593] + MEM[8594];
assign MEM[8690] = MEM[8624] + MEM[8625];
assign MEM[8691] = MEM[8628] + MEM[8629];
assign MEM[8692] = MEM[8634] + MEM[8635];
assign MEM[8693] = MEM[8680] + MEM[7259];
assign MEM[8694] = MEM[45] + MEM[3847];
assign MEM[8695] = MEM[54] + MEM[600];
assign MEM[8696] = MEM[63] + MEM[3858];
assign MEM[8697] = MEM[79] + MEM[1774];
assign MEM[8698] = MEM[87] + MEM[2462];
assign MEM[8699] = MEM[127] + MEM[4061];
assign MEM[8700] = MEM[134] + MEM[4782];
assign MEM[8701] = MEM[136] + MEM[137];
assign MEM[8702] = MEM[138] + MEM[139];
assign MEM[8703] = MEM[140] + MEM[8701];
assign MEM[8704] = MEM[151] + MEM[3335];
assign MEM[8705] = MEM[182] + MEM[1166];
assign MEM[8706] = MEM[295] + MEM[4414];
assign MEM[8707] = MEM[315] + MEM[3309];
assign MEM[8708] = MEM[318] + MEM[395];
assign MEM[8709] = MEM[323] + MEM[1283];
assign MEM[8710] = MEM[357] + MEM[3357];
assign MEM[8711] = MEM[380] + MEM[5109];
assign MEM[8712] = MEM[412] + MEM[4238];
assign MEM[8713] = MEM[526] + MEM[709];
assign MEM[8714] = MEM[601] + MEM[2323];
assign MEM[8715] = MEM[602] + MEM[3476];
assign MEM[8716] = MEM[620] + MEM[1195];
assign MEM[8717] = MEM[655] + MEM[3397];
assign MEM[8718] = MEM[782] + MEM[3874];
assign MEM[8719] = MEM[805] + MEM[4653];
assign MEM[8720] = MEM[887] + MEM[4798];
assign MEM[8721] = MEM[1012] + MEM[2958];
assign MEM[8722] = MEM[1015] + MEM[3239];
assign MEM[8723] = MEM[1018] + MEM[5779];
assign MEM[8724] = MEM[1023] + MEM[1687];
assign MEM[8725] = MEM[1029] + MEM[1486];
assign MEM[8726] = MEM[1063] + MEM[5928];
assign MEM[8727] = MEM[1101] + MEM[4202];
assign MEM[8728] = MEM[1151] + MEM[5694];
assign MEM[8729] = MEM[1203] + MEM[327];
assign MEM[8730] = MEM[1221] + MEM[1998];
assign MEM[8731] = MEM[1270] + MEM[3614];
assign MEM[8732] = MEM[1317] + MEM[5937];
assign MEM[8733] = MEM[1320] + MEM[1321];
assign MEM[8734] = MEM[1323] + MEM[2605];
assign MEM[8735] = MEM[1334] + MEM[2797];
assign MEM[8736] = MEM[1375] + MEM[1603];
assign MEM[8737] = MEM[1436] + MEM[3340];
assign MEM[8738] = MEM[1453] + MEM[3199];
assign MEM[8739] = MEM[1469] + MEM[2125];
assign MEM[8740] = MEM[1500] + MEM[6556];
assign MEM[8741] = MEM[1522] + MEM[1618];
assign MEM[8742] = MEM[1538] + MEM[5075];
assign MEM[8743] = MEM[1554] + MEM[958];
assign MEM[8744] = MEM[1587] + MEM[2946];
assign MEM[8745] = MEM[1631] + MEM[3963];
assign MEM[8746] = MEM[1658] + MEM[8226];
assign MEM[8747] = MEM[1707] + MEM[3010];
assign MEM[8748] = MEM[1743] + MEM[2140];
assign MEM[8749] = MEM[1751] + MEM[3341];
assign MEM[8750] = MEM[1764] + MEM[3093];
assign MEM[8751] = MEM[1766] + MEM[5847];
assign MEM[8752] = MEM[1773] + MEM[5511];
assign MEM[8753] = MEM[1799] + MEM[3210];
assign MEM[8754] = MEM[1803] + MEM[5973];
assign MEM[8755] = MEM[1860] + MEM[2999];
assign MEM[8756] = MEM[1870] + MEM[6629];
assign MEM[8757] = MEM[1907] + MEM[403];
assign MEM[8758] = MEM[1934] + MEM[2004];
assign MEM[8759] = MEM[1942] + MEM[4901];
assign MEM[8760] = MEM[1950] + MEM[5222];
assign MEM[8761] = MEM[1997] + MEM[6205];
assign MEM[8762] = MEM[2052] + MEM[2198];
assign MEM[8763] = MEM[2107] + MEM[2819];
assign MEM[8764] = MEM[2115] + MEM[4214];
assign MEM[8765] = MEM[2117] + MEM[2453];
assign MEM[8766] = MEM[2180] + MEM[4574];
assign MEM[8767] = MEM[2205] + MEM[2510];
assign MEM[8768] = MEM[2214] + MEM[3163];
assign MEM[8769] = MEM[2308] + MEM[754];
assign MEM[8770] = MEM[2310] + MEM[2550];
assign MEM[8771] = MEM[2316] + MEM[4157];
assign MEM[8772] = MEM[2335] + MEM[3298];
assign MEM[8773] = MEM[2434] + MEM[4650];
assign MEM[8774] = MEM[2485] + MEM[4246];
assign MEM[8775] = MEM[2494] + MEM[3879];
assign MEM[8776] = MEM[2522] + MEM[2523];
assign MEM[8777] = MEM[2524] + MEM[6569];
assign MEM[8778] = MEM[2540] + MEM[4180];
assign MEM[8779] = MEM[2567] + MEM[4764];
assign MEM[8780] = MEM[2580] + MEM[2245];
assign MEM[8781] = MEM[2590] + MEM[5348];
assign MEM[8782] = MEM[2611] + MEM[3275];
assign MEM[8783] = MEM[2676] + MEM[3111];
assign MEM[8784] = MEM[2732] + MEM[3279];
assign MEM[8785] = MEM[2740] + MEM[5354];
assign MEM[8786] = MEM[2783] + MEM[5654];
assign MEM[8787] = MEM[2822] + MEM[4702];
assign MEM[8788] = MEM[2834] + MEM[2835];
assign MEM[8789] = MEM[2837] + MEM[2820];
assign MEM[8790] = MEM[2839] + MEM[1206];
assign MEM[8791] = MEM[2866] + MEM[2876];
assign MEM[8792] = MEM[2870] + MEM[6613];
assign MEM[8793] = MEM[2887] + MEM[5015];
assign MEM[8794] = MEM[2895] + MEM[2930];
assign MEM[8795] = MEM[2900] + MEM[5102];
assign MEM[8796] = MEM[2933] + MEM[5246];
assign MEM[8797] = MEM[2950] + MEM[6007];
assign MEM[8798] = MEM[3020] + MEM[6037];
assign MEM[8799] = MEM[3030] + MEM[6812];
assign MEM[8800] = MEM[3109] + MEM[5356];
assign MEM[8801] = MEM[3189] + MEM[3259];
assign MEM[8802] = MEM[3308] + MEM[5930];
assign MEM[8803] = MEM[3324] + MEM[4522];
assign MEM[8804] = MEM[3327] + MEM[3230];
assign MEM[8805] = MEM[3347] + MEM[2350];
assign MEM[8806] = MEM[3358] + MEM[6149];
assign MEM[8807] = MEM[3415] + MEM[5509];
assign MEM[8808] = MEM[3419] + MEM[3418];
assign MEM[8809] = MEM[3483] + MEM[3482];
assign MEM[8810] = MEM[3547] + MEM[5405];
assign MEM[8811] = MEM[3670] + MEM[5695];
assign MEM[8812] = MEM[3757] + MEM[4486];
assign MEM[8813] = MEM[3816] + MEM[3817];
assign MEM[8814] = MEM[3818] + MEM[3819];
assign MEM[8815] = MEM[3820] + MEM[8813];
assign MEM[8816] = MEM[3850] + MEM[6738];
assign MEM[8817] = MEM[3854] + MEM[837];
assign MEM[8818] = MEM[3866] + MEM[6586];
assign MEM[8819] = MEM[3927] + MEM[5051];
assign MEM[8820] = MEM[3930] + MEM[1989];
assign MEM[8821] = MEM[3936] + MEM[3937];
assign MEM[8822] = MEM[3967] + MEM[818];
assign MEM[8823] = MEM[3999] + MEM[5115];
assign MEM[8824] = MEM[4020] + MEM[973];
assign MEM[8825] = MEM[4040] + MEM[4041];
assign MEM[8826] = MEM[4042] + MEM[4043];
assign MEM[8827] = MEM[4053] + MEM[1388];
assign MEM[8828] = MEM[4076] + MEM[5122];
assign MEM[8829] = MEM[4141] + MEM[3654];
assign MEM[8830] = MEM[4142] + MEM[5670];
assign MEM[8831] = MEM[4179] + MEM[7250];
assign MEM[8832] = MEM[4253] + MEM[1187];
assign MEM[8833] = MEM[4255] + MEM[5084];
assign MEM[8834] = MEM[4301] + MEM[4676];
assign MEM[8835] = MEM[4311] + MEM[6179];
assign MEM[8836] = MEM[4322] + MEM[5557];
assign MEM[8837] = MEM[4324] + MEM[3150];
assign MEM[8838] = MEM[4326] + MEM[142];
assign MEM[8839] = MEM[4371] + MEM[4386];
assign MEM[8840] = MEM[4395] + MEM[4394];
assign MEM[8841] = MEM[4405] + MEM[5735];
assign MEM[8842] = MEM[4470] + MEM[4501];
assign MEM[8843] = MEM[4490] + MEM[4884];
assign MEM[8844] = MEM[4507] + MEM[4669];
assign MEM[8845] = MEM[4508] + MEM[6659];
assign MEM[8846] = MEM[4659] + MEM[1678];
assign MEM[8847] = MEM[4703] + MEM[2206];
assign MEM[8848] = MEM[4748] + MEM[951];
assign MEM[8849] = MEM[4749] + MEM[3723];
assign MEM[8850] = MEM[4771] + MEM[1750];
assign MEM[8851] = MEM[4836] + MEM[1662];
assign MEM[8852] = MEM[4867] + MEM[3268];
assign MEM[8853] = MEM[4934] + MEM[5875];
assign MEM[8854] = MEM[4978] + MEM[5914];
assign MEM[8855] = MEM[5008] + MEM[5009];
assign MEM[8856] = MEM[5014] + MEM[5053];
assign MEM[8857] = MEM[5062] + MEM[6237];
assign MEM[8858] = MEM[5092] + MEM[5415];
assign MEM[8859] = MEM[5093] + MEM[6223];
assign MEM[8860] = MEM[5119] + MEM[3310];
assign MEM[8861] = MEM[5172] + MEM[6609];
assign MEM[8862] = MEM[5174] + MEM[3901];
assign MEM[8863] = MEM[5223] + MEM[4691];
assign MEM[8864] = MEM[5262] + MEM[6061];
assign MEM[8865] = MEM[5309] + MEM[6614];
assign MEM[8866] = MEM[5347] + MEM[2191];
assign MEM[8867] = MEM[5376] + MEM[5377];
assign MEM[8868] = MEM[5378] + MEM[5379];
assign MEM[8869] = MEM[5380] + MEM[8867];
assign MEM[8870] = MEM[5420] + MEM[1605];
assign MEM[8871] = MEM[5475] + MEM[1535];
assign MEM[8872] = MEM[5494] + MEM[1946];
assign MEM[8873] = MEM[5562] + MEM[3613];
assign MEM[8874] = MEM[5614] + MEM[3523];
assign MEM[8875] = MEM[5630] + MEM[2131];
assign MEM[8876] = MEM[5650] + MEM[4717];
assign MEM[8877] = MEM[5660] + MEM[1292];
assign MEM[8878] = MEM[5661] + MEM[787];
assign MEM[8879] = MEM[5699] + MEM[1735];
assign MEM[8880] = MEM[5701] + MEM[3911];
assign MEM[8881] = MEM[5750] + MEM[5331];
assign MEM[8882] = MEM[5821] + MEM[7071];
assign MEM[8883] = MEM[5845] + MEM[1879];
assign MEM[8884] = MEM[5854] + MEM[1186];
assign MEM[8885] = MEM[5868] + MEM[5252];
assign MEM[8886] = MEM[5904] + MEM[1987];
assign MEM[8887] = MEM[5933] + MEM[2139];
assign MEM[8888] = MEM[5935] + MEM[6961];
assign MEM[8889] = MEM[5957] + MEM[3293];
assign MEM[8890] = MEM[5970] + MEM[469];
assign MEM[8891] = MEM[5971] + MEM[2534];
assign MEM[8892] = MEM[6011] + MEM[6188];
assign MEM[8893] = MEM[6024] + MEM[6025];
assign MEM[8894] = MEM[6026] + MEM[6027];
assign MEM[8895] = MEM[6028] + MEM[8893];
assign MEM[8896] = MEM[6093] + MEM[6206];
assign MEM[8897] = MEM[6117] + MEM[6912];
assign MEM[8898] = MEM[6130] + MEM[1326];
assign MEM[8899] = MEM[6164] + MEM[6198];
assign MEM[8900] = MEM[6190] + MEM[4462];
assign MEM[8901] = MEM[6519] + MEM[2988];
assign MEM[8902] = MEM[6560] + MEM[1902];
assign MEM[8903] = MEM[6561] + MEM[6693];
assign MEM[8904] = MEM[6568] + MEM[158];
assign MEM[8905] = MEM[6579] + MEM[1756];
assign MEM[8906] = MEM[6610] + MEM[3668];
assign MEM[8907] = MEM[6611] + MEM[2426];
assign MEM[8908] = MEM[6615] + MEM[2164];
assign MEM[8909] = MEM[6617] + MEM[285];
assign MEM[8910] = MEM[6619] + MEM[6697];
assign MEM[8911] = MEM[6633] + MEM[6871];
assign MEM[8912] = MEM[6635] + MEM[2558];
assign MEM[8913] = MEM[6648] + MEM[6842];
assign MEM[8914] = MEM[6660] + MEM[4124];
assign MEM[8915] = MEM[6674] + MEM[1580];
assign MEM[8916] = MEM[6677] + MEM[4181];
assign MEM[8917] = MEM[6678] + MEM[6828];
assign MEM[8918] = MEM[6685] + MEM[5230];
assign MEM[8919] = MEM[6701] + MEM[5693];
assign MEM[8920] = MEM[6705] + MEM[7016];
assign MEM[8921] = MEM[6707] + MEM[7160];
assign MEM[8922] = MEM[6710] + MEM[4979];
assign MEM[8923] = MEM[6736] + MEM[3543];
assign MEM[8924] = MEM[6748] + MEM[6992];
assign MEM[8925] = MEM[6752] + MEM[4389];
assign MEM[8926] = MEM[6776] + MEM[6929];
assign MEM[8927] = MEM[6796] + MEM[3710];
assign MEM[8928] = MEM[6799] + MEM[6939];
assign MEM[8929] = MEM[6809] + MEM[5364];
assign MEM[8930] = MEM[6817] + MEM[6880];
assign MEM[8931] = MEM[6827] + MEM[6831];
assign MEM[8932] = MEM[6840] + MEM[6839];
assign MEM[8933] = MEM[6845] + MEM[29];
assign MEM[8934] = MEM[6847] + MEM[4223];
assign MEM[8935] = MEM[6866] + MEM[4722];
assign MEM[8936] = MEM[6872] + MEM[7005];
assign MEM[8937] = MEM[6874] + MEM[5098];
assign MEM[8938] = MEM[6885] + MEM[2087];
assign MEM[8939] = MEM[6889] + MEM[6836];
assign MEM[8940] = MEM[6899] + MEM[7379];
assign MEM[8941] = MEM[6911] + MEM[271];
assign MEM[8942] = MEM[6932] + MEM[585];
assign MEM[8943] = MEM[6933] + MEM[6931];
assign MEM[8944] = MEM[6950] + MEM[6656];
assign MEM[8945] = MEM[6955] + MEM[2647];
assign MEM[8946] = MEM[6971] + MEM[2218];
assign MEM[8947] = MEM[6982] + MEM[7125];
assign MEM[8948] = MEM[6997] + MEM[6675];
assign MEM[8949] = MEM[7041] + MEM[7356];
assign MEM[8950] = MEM[7070] + MEM[722];
assign MEM[8951] = MEM[7233] + MEM[6741];
assign MEM[8952] = MEM[7255] + MEM[1602];
assign MEM[8953] = MEM[8702] + MEM[8703];
assign MEM[8954] = MEM[8776] + MEM[7117];
assign MEM[8955] = MEM[8794] + MEM[6826];
assign MEM[8956] = MEM[8809] + MEM[7506];
assign MEM[8957] = MEM[8814] + MEM[8815];
assign MEM[8958] = MEM[8825] + MEM[8826];
assign MEM[8959] = MEM[8840] + MEM[7533];
assign MEM[8960] = MEM[8855] + MEM[5010];
assign MEM[8961] = MEM[8868] + MEM[8869];
assign MEM[8962] = MEM[8894] + MEM[8895];
assign MEM[8963] = MEM[21] + MEM[2722];
assign MEM[8964] = MEM[48] + MEM[49];
assign MEM[8965] = MEM[50] + MEM[51];
assign MEM[8966] = MEM[52] + MEM[8964];
assign MEM[8967] = MEM[107] + MEM[885];
assign MEM[8968] = MEM[116] + MEM[5111];
assign MEM[8969] = MEM[150] + MEM[5351];
assign MEM[8970] = MEM[174] + MEM[4495];
assign MEM[8971] = MEM[190] + MEM[283];
assign MEM[8972] = MEM[239] + MEM[1780];
assign MEM[8973] = MEM[263] + MEM[5202];
assign MEM[8974] = MEM[277] + MEM[5469];
assign MEM[8975] = MEM[293] + MEM[3118];
assign MEM[8976] = MEM[324] + MEM[583];
assign MEM[8977] = MEM[351] + MEM[2166];
assign MEM[8978] = MEM[364] + MEM[5519];
assign MEM[8979] = MEM[388] + MEM[1260];
assign MEM[8980] = MEM[518] + MEM[5955];
assign MEM[8981] = MEM[572] + MEM[3054];
assign MEM[8982] = MEM[610] + MEM[1591];
assign MEM[8983] = MEM[639] + MEM[2378];
assign MEM[8984] = MEM[669] + MEM[2266];
assign MEM[8985] = MEM[747] + MEM[5471];
assign MEM[8986] = MEM[773] + MEM[2869];
assign MEM[8987] = MEM[790] + MEM[4572];
assign MEM[8988] = MEM[829] + MEM[3092];
assign MEM[8989] = MEM[834] + MEM[5773];
assign MEM[8990] = MEM[845] + MEM[5506];
assign MEM[8991] = MEM[910] + MEM[1957];
assign MEM[8992] = MEM[947] + MEM[1300];
assign MEM[8993] = MEM[987] + MEM[2246];
assign MEM[8994] = MEM[988] + MEM[1450];
assign MEM[8995] = MEM[1034] + MEM[2444];
assign MEM[8996] = MEM[1044] + MEM[4742];
assign MEM[8997] = MEM[1059] + MEM[3583];
assign MEM[8998] = MEM[1084] + MEM[2044];
assign MEM[8999] = MEM[1181] + MEM[3318];
assign MEM[9000] = MEM[1198] + MEM[1382];
assign MEM[9001] = MEM[1205] + MEM[3605];
assign MEM[9002] = MEM[1231] + MEM[2942];
assign MEM[9003] = MEM[1234] + MEM[1235];
assign MEM[9004] = MEM[1276] + MEM[1567];
assign MEM[9005] = MEM[1294] + MEM[1309];
assign MEM[9006] = MEM[1342] + MEM[2326];
assign MEM[9007] = MEM[1378] + MEM[6062];
assign MEM[9008] = MEM[1397] + MEM[2358];
assign MEM[9009] = MEM[1398] + MEM[4175];
assign MEM[9010] = MEM[1410] + MEM[5795];
assign MEM[9011] = MEM[1423] + MEM[4055];
assign MEM[9012] = MEM[1437] + MEM[4741];
assign MEM[9013] = MEM[1451] + MEM[3799];
assign MEM[9014] = MEM[1503] + MEM[4891];
assign MEM[9015] = MEM[1517] + MEM[4950];
assign MEM[9016] = MEM[1519] + MEM[5446];
assign MEM[9017] = MEM[1526] + MEM[2318];
assign MEM[9018] = MEM[1628] + MEM[4196];
assign MEM[9019] = MEM[1650] + MEM[2045];
assign MEM[9020] = MEM[1659] + MEM[2903];
assign MEM[9021] = MEM[1717] + MEM[2621];
assign MEM[9022] = MEM[1723] + MEM[2549];
assign MEM[9023] = MEM[1727] + MEM[199];
assign MEM[9024] = MEM[1778] + MEM[5908];
assign MEM[9025] = MEM[1828] + MEM[6012];
assign MEM[9026] = MEM[1830] + MEM[5710];
assign MEM[9027] = MEM[1852] + MEM[3437];
assign MEM[9028] = MEM[1892] + MEM[5023];
assign MEM[9029] = MEM[1967] + MEM[2239];
assign MEM[9030] = MEM[1982] + MEM[5983];
assign MEM[9031] = MEM[1995] + MEM[5207];
assign MEM[9032] = MEM[2031] + MEM[3299];
assign MEM[9033] = MEM[2078] + MEM[6745];
assign MEM[9034] = MEM[2084] + MEM[5772];
assign MEM[9035] = MEM[2095] + MEM[5389];
assign MEM[9036] = MEM[2101] + MEM[3471];
assign MEM[9037] = MEM[2181] + MEM[2491];
assign MEM[9038] = MEM[2199] + MEM[2406];
assign MEM[9039] = MEM[2226] + MEM[4278];
assign MEM[9040] = MEM[2290] + MEM[2291];
assign MEM[9041] = MEM[2306] + MEM[4970];
assign MEM[9042] = MEM[2314] + MEM[3781];
assign MEM[9043] = MEM[2338] + MEM[3679];
assign MEM[9044] = MEM[2359] + MEM[4071];
assign MEM[9045] = MEM[2375] + MEM[4796];
assign MEM[9046] = MEM[2380] + MEM[2430];
assign MEM[9047] = MEM[2381] + MEM[5886];
assign MEM[9048] = MEM[2390] + MEM[2931];
assign MEM[9049] = MEM[2399] + MEM[2830];
assign MEM[9050] = MEM[2431] + MEM[6558];
assign MEM[9051] = MEM[2459] + MEM[6022];
assign MEM[9052] = MEM[2471] + MEM[3108];
assign MEM[9053] = MEM[2477] + MEM[4091];
assign MEM[9054] = MEM[2495] + MEM[2766];
assign MEM[9055] = MEM[2506] + MEM[2702];
assign MEM[9056] = MEM[2508] + MEM[4511];
assign MEM[9057] = MEM[2573] + MEM[6749];
assign MEM[9058] = MEM[2588] + MEM[6620];
assign MEM[9059] = MEM[2723] + MEM[2862];
assign MEM[9060] = MEM[2735] + MEM[4468];
assign MEM[9061] = MEM[2743] + MEM[6700];
assign MEM[9062] = MEM[2751] + MEM[1806];
assign MEM[9063] = MEM[2846] + MEM[4340];
assign MEM[9064] = MEM[2891] + MEM[2037];
assign MEM[9065] = MEM[2894] + MEM[5414];
assign MEM[9066] = MEM[2934] + MEM[5213];
assign MEM[9067] = MEM[3039] + MEM[6751];
assign MEM[9068] = MEM[3094] + MEM[6698];
assign MEM[9069] = MEM[3114] + MEM[3714];
assign MEM[9070] = MEM[3179] + MEM[5675];
assign MEM[9071] = MEM[3194] + MEM[6709];
assign MEM[9072] = MEM[3247] + MEM[2483];
assign MEM[9073] = MEM[3262] + MEM[4461];
assign MEM[9074] = MEM[3284] + MEM[3764];
assign MEM[9075] = MEM[3342] + MEM[6532];
assign MEM[9076] = MEM[3351] + MEM[4460];
assign MEM[9077] = MEM[3374] + MEM[5006];
assign MEM[9078] = MEM[3380] + MEM[4101];
assign MEM[9079] = MEM[3394] + MEM[927];
assign MEM[9080] = MEM[3422] + MEM[5929];
assign MEM[9081] = MEM[3427] + MEM[6085];
assign MEM[9082] = MEM[3435] + MEM[2726];
assign MEM[9083] = MEM[3452] + MEM[6715];
assign MEM[9084] = MEM[3458] + MEM[5244];
assign MEM[9085] = MEM[3479] + MEM[3095];
assign MEM[9086] = MEM[3486] + MEM[4687];
assign MEM[9087] = MEM[3500] + MEM[2050];
assign MEM[9088] = MEM[3503] + MEM[247];
assign MEM[9089] = MEM[3533] + MEM[5739];
assign MEM[9090] = MEM[3539] + MEM[4862];
assign MEM[9091] = MEM[3581] + MEM[5086];
assign MEM[9092] = MEM[3631] + MEM[6229];
assign MEM[9093] = MEM[3634] + MEM[2811];
assign MEM[9094] = MEM[3650] + MEM[4341];
assign MEM[9095] = MEM[3660] + MEM[39];
assign MEM[9096] = MEM[3671] + MEM[6172];
assign MEM[9097] = MEM[3692] + MEM[4295];
assign MEM[9098] = MEM[3724] + MEM[5756];
assign MEM[9099] = MEM[3726] + MEM[3990];
assign MEM[9100] = MEM[3766] + MEM[3261];
assign MEM[9101] = MEM[3770] + MEM[5678];
assign MEM[9102] = MEM[3780] + MEM[2006];
assign MEM[9103] = MEM[3868] + MEM[4243];
assign MEM[9104] = MEM[3938] + MEM[8821];
assign MEM[9105] = MEM[3974] + MEM[6717];
assign MEM[9106] = MEM[3991] + MEM[4629];
assign MEM[9107] = MEM[4021] + MEM[694];
assign MEM[9108] = MEM[4067] + MEM[5903];
assign MEM[9109] = MEM[4077] + MEM[5100];
assign MEM[9110] = MEM[4131] + MEM[5306];
assign MEM[9111] = MEM[4212] + MEM[6900];
assign MEM[9112] = MEM[4215] + MEM[3084];
assign MEM[9113] = MEM[4268] + MEM[4347];
assign MEM[9114] = MEM[4358] + MEM[1565];
assign MEM[9115] = MEM[4382] + MEM[2586];
assign MEM[9116] = MEM[4423] + MEM[6046];
assign MEM[9117] = MEM[4454] + MEM[303];
assign MEM[9118] = MEM[4549] + MEM[2396];
assign MEM[9119] = MEM[4567] + MEM[2438];
assign MEM[9120] = MEM[4575] + MEM[5131];
assign MEM[9121] = MEM[4695] + MEM[2578];
assign MEM[9122] = MEM[4715] + MEM[5539];
assign MEM[9123] = MEM[4727] + MEM[786];
assign MEM[9124] = MEM[4740] + MEM[5495];
assign MEM[9125] = MEM[4751] + MEM[7286];
assign MEM[9126] = MEM[4767] + MEM[5106];
assign MEM[9127] = MEM[4786] + MEM[4900];
assign MEM[9128] = MEM[4831] + MEM[3783];
assign MEM[9129] = MEM[4859] + MEM[4858];
assign MEM[9130] = MEM[4869] + MEM[3119];
assign MEM[9131] = MEM[4886] + MEM[4434];
assign MEM[9132] = MEM[4982] + MEM[2330];
assign MEM[9133] = MEM[4988] + MEM[5476];
assign MEM[9134] = MEM[5004] + MEM[6101];
assign MEM[9135] = MEM[5016] + MEM[5017];
assign MEM[9136] = MEM[5027] + MEM[1627];
assign MEM[9137] = MEM[5085] + MEM[1109];
assign MEM[9138] = MEM[5125] + MEM[3959];
assign MEM[9139] = MEM[5190] + MEM[4125];
assign MEM[9140] = MEM[5191] + MEM[6905];
assign MEM[9141] = MEM[5295] + MEM[7170];
assign MEM[9142] = MEM[5316] + MEM[742];
assign MEM[9143] = MEM[5442] + MEM[4965];
assign MEM[9144] = MEM[5499] + MEM[844];
assign MEM[9145] = MEM[5518] + MEM[1970];
assign MEM[9146] = MEM[5531] + MEM[6652];
assign MEM[9147] = MEM[5551] + MEM[4949];
assign MEM[9148] = MEM[5567] + MEM[5703];
assign MEM[9149] = MEM[5571] + MEM[6087];
assign MEM[9150] = MEM[5615] + MEM[1663];
assign MEM[9151] = MEM[5651] + MEM[3563];
assign MEM[9152] = MEM[5813] + MEM[2599];
assign MEM[9153] = MEM[5869] + MEM[4146];
assign MEM[9154] = MEM[5905] + MEM[5906];
assign MEM[9155] = MEM[5917] + MEM[4879];
assign MEM[9156] = MEM[5959] + MEM[6916];
assign MEM[9157] = MEM[5962] + MEM[7058];
assign MEM[9158] = MEM[5974] + MEM[1022];
assign MEM[9159] = MEM[5989] + MEM[3069];
assign MEM[9160] = MEM[6003] + MEM[1108];
assign MEM[9161] = MEM[6077] + MEM[1222];
assign MEM[9162] = MEM[6080] + MEM[6081];
assign MEM[9163] = MEM[6082] + MEM[6083];
assign MEM[9164] = MEM[6084] + MEM[9162];
assign MEM[9165] = MEM[6131] + MEM[6816];
assign MEM[9166] = MEM[6151] + MEM[6170];
assign MEM[9167] = MEM[6187] + MEM[4494];
assign MEM[9168] = MEM[6191] + MEM[2331];
assign MEM[9169] = MEM[6518] + MEM[404];
assign MEM[9170] = MEM[6616] + MEM[5290];
assign MEM[9171] = MEM[6644] + MEM[875];
assign MEM[9172] = MEM[6649] + MEM[1623];
assign MEM[9173] = MEM[6658] + MEM[4133];
assign MEM[9174] = MEM[6670] + MEM[5300];
assign MEM[9175] = MEM[6681] + MEM[3739];
assign MEM[9176] = MEM[6682] + MEM[3269];
assign MEM[9177] = MEM[6691] + MEM[851];
assign MEM[9178] = MEM[6703] + MEM[6744];
assign MEM[9179] = MEM[6706] + MEM[4607];
assign MEM[9180] = MEM[6714] + MEM[2884];
assign MEM[9181] = MEM[6718] + MEM[2731];
assign MEM[9182] = MEM[6725] + MEM[6886];
assign MEM[9183] = MEM[6729] + MEM[6740];
assign MEM[9184] = MEM[6743] + MEM[613];
assign MEM[9185] = MEM[6753] + MEM[4535];
assign MEM[9186] = MEM[6754] + MEM[4194];
assign MEM[9187] = MEM[6787] + MEM[6848];
assign MEM[9188] = MEM[6795] + MEM[6804];
assign MEM[9189] = MEM[6813] + MEM[2514];
assign MEM[9190] = MEM[6814] + MEM[2813];
assign MEM[9191] = MEM[6819] + MEM[5486];
assign MEM[9192] = MEM[6837] + MEM[2220];
assign MEM[9193] = MEM[6858] + MEM[3174];
assign MEM[9194] = MEM[6859] + MEM[2167];
assign MEM[9195] = MEM[6887] + MEM[6775];
assign MEM[9196] = MEM[6898] + MEM[3540];
assign MEM[9197] = MEM[6903] + MEM[2669];
assign MEM[9198] = MEM[6910] + MEM[2964];
assign MEM[9199] = MEM[6917] + MEM[5927];
assign MEM[9200] = MEM[6940] + MEM[7184];
assign MEM[9201] = MEM[6943] + MEM[6952];
assign MEM[9202] = MEM[6944] + MEM[1259];
assign MEM[9203] = MEM[6958] + MEM[5255];
assign MEM[9204] = MEM[6962] + MEM[341];
assign MEM[9205] = MEM[6970] + MEM[4147];
assign MEM[9206] = MEM[6986] + MEM[3203];
assign MEM[9207] = MEM[6987] + MEM[2901];
assign MEM[9208] = MEM[7002] + MEM[4898];
assign MEM[9209] = MEM[7018] + MEM[6086];
assign MEM[9210] = MEM[7022] + MEM[3423];
assign MEM[9211] = MEM[7049] + MEM[7056];
assign MEM[9212] = MEM[7050] + MEM[7522];
assign MEM[9213] = MEM[7069] + MEM[4516];
assign MEM[9214] = MEM[7089] + MEM[5266];
assign MEM[9215] = MEM[7202] + MEM[5383];
assign MEM[9216] = MEM[7203] + MEM[7040];
assign MEM[9217] = MEM[7258] + MEM[7449];
assign MEM[9218] = MEM[7445] + MEM[6849];
assign MEM[9219] = MEM[8965] + MEM[8966];
assign MEM[9220] = MEM[9040] + MEM[7274];
assign MEM[9221] = MEM[9135] + MEM[5018];
assign MEM[9222] = MEM[9163] + MEM[9164];
assign MEM[9223] = MEM[5] + MEM[262];
assign MEM[9224] = MEM[22] + MEM[423];
assign MEM[9225] = MEM[64] + MEM[65];
assign MEM[9226] = MEM[66] + MEM[67];
assign MEM[9227] = MEM[68] + MEM[9225];
assign MEM[9228] = MEM[70] + MEM[803];
assign MEM[9229] = MEM[118] + MEM[2883];
assign MEM[9230] = MEM[215] + MEM[3028];
assign MEM[9231] = MEM[245] + MEM[2618];
assign MEM[9232] = MEM[279] + MEM[878];
assign MEM[9233] = MEM[309] + MEM[4822];
assign MEM[9234] = MEM[399] + MEM[2603];
assign MEM[9235] = MEM[405] + MEM[3557];
assign MEM[9236] = MEM[454] + MEM[6661];
assign MEM[9237] = MEM[522] + MEM[7141];
assign MEM[9238] = MEM[538] + MEM[6755];
assign MEM[9239] = MEM[541] + MEM[2268];
assign MEM[9240] = MEM[580] + MEM[2270];
assign MEM[9241] = MEM[594] + MEM[1275];
assign MEM[9242] = MEM[701] + MEM[3877];
assign MEM[9243] = MEM[743] + MEM[1583];
assign MEM[9244] = MEM[756] + MEM[1413];
assign MEM[9245] = MEM[794] + MEM[2484];
assign MEM[9246] = MEM[799] + MEM[1677];
assign MEM[9247] = MEM[813] + MEM[2317];
assign MEM[9248] = MEM[838] + MEM[1741];
assign MEM[9249] = MEM[866] + MEM[6747];
assign MEM[9250] = MEM[867] + MEM[3302];
assign MEM[9251] = MEM[918] + MEM[6746];
assign MEM[9252] = MEM[940] + MEM[5770];
assign MEM[9253] = MEM[950] + MEM[5980];
assign MEM[9254] = MEM[1005] + MEM[4204];
assign MEM[9255] = MEM[1011] + MEM[2414];
assign MEM[9256] = MEM[1019] + MEM[2476];
assign MEM[9257] = MEM[1027] + MEM[2627];
assign MEM[9258] = MEM[1070] + MEM[2878];
assign MEM[9259] = MEM[1071] + MEM[4149];
assign MEM[9260] = MEM[1076] + MEM[3698];
assign MEM[9261] = MEM[1095] + MEM[5037];
assign MEM[9262] = MEM[1183] + MEM[6808];
assign MEM[9263] = MEM[1215] + MEM[5831];
assign MEM[9264] = MEM[1219] + MEM[5335];
assign MEM[9265] = MEM[1247] + MEM[1351];
assign MEM[9266] = MEM[1262] + MEM[3926];
assign MEM[9267] = MEM[1363] + MEM[2173];
assign MEM[9268] = MEM[1462] + MEM[3510];
assign MEM[9269] = MEM[1508] + MEM[2030];
assign MEM[9270] = MEM[1548] + MEM[3651];
assign MEM[9271] = MEM[1613] + MEM[5291];
assign MEM[9272] = MEM[1642] + MEM[7132];
assign MEM[9273] = MEM[1702] + MEM[2845];
assign MEM[9274] = MEM[1746] + MEM[3323];
assign MEM[9275] = MEM[1757] + MEM[3185];
assign MEM[9276] = MEM[1782] + MEM[4189];
assign MEM[9277] = MEM[1813] + MEM[2038];
assign MEM[9278] = MEM[1819] + MEM[4316];
assign MEM[9279] = MEM[1846] + MEM[7012];
assign MEM[9280] = MEM[1917] + MEM[5437];
assign MEM[9281] = MEM[1924] + MEM[4957];
assign MEM[9282] = MEM[1947] + MEM[1754];
assign MEM[9283] = MEM[1962] + MEM[2186];
assign MEM[9284] = MEM[1966] + MEM[2299];
assign MEM[9285] = MEM[2100] + MEM[5423];
assign MEM[9286] = MEM[2174] + MEM[3285];
assign MEM[9287] = MEM[2183] + MEM[2677];
assign MEM[9288] = MEM[2187] + MEM[4802];
assign MEM[9289] = MEM[2196] + MEM[2788];
assign MEM[9290] = MEM[2219] + MEM[6271];
assign MEM[9291] = MEM[2230] + MEM[6942];
assign MEM[9292] = MEM[2237] + MEM[6875];
assign MEM[9293] = MEM[2260] + MEM[5332];
assign MEM[9294] = MEM[2261] + MEM[5396];
assign MEM[9295] = MEM[2262] + MEM[5117];
assign MEM[9296] = MEM[2274] + MEM[5736];
assign MEM[9297] = MEM[2364] + MEM[5116];
assign MEM[9298] = MEM[2366] + MEM[5683];
assign MEM[9299] = MEM[2394] + MEM[1684];
assign MEM[9300] = MEM[2436] + MEM[1179];
assign MEM[9301] = MEM[2451] + MEM[5043];
assign MEM[9302] = MEM[2517] + MEM[5118];
assign MEM[9303] = MEM[2575] + MEM[3546];
assign MEM[9304] = MEM[2581] + MEM[607];
assign MEM[9305] = MEM[2589] + MEM[3243];
assign MEM[9306] = MEM[2631] + MEM[1372];
assign MEM[9307] = MEM[2668] + MEM[5087];
assign MEM[9308] = MEM[2684] + MEM[5254];
assign MEM[9309] = MEM[2741] + MEM[6888];
assign MEM[9310] = MEM[2802] + MEM[3127];
assign MEM[9311] = MEM[2803] + MEM[6857];
assign MEM[9312] = MEM[2810] + MEM[5175];
assign MEM[9313] = MEM[2826] + MEM[2827];
assign MEM[9314] = MEM[2838] + MEM[3278];
assign MEM[9315] = MEM[2935] + MEM[4244];
assign MEM[9316] = MEM[2941] + MEM[7193];
assign MEM[9317] = MEM[2970] + MEM[7035];
assign MEM[9318] = MEM[3018] + MEM[6981];
assign MEM[9319] = MEM[3035] + MEM[6921];
assign MEM[9320] = MEM[3037] + MEM[1148];
assign MEM[9321] = MEM[3055] + MEM[3143];
assign MEM[9322] = MEM[3106] + MEM[3915];
assign MEM[9323] = MEM[3171] + MEM[3519];
assign MEM[9324] = MEM[3180] + MEM[3372];
assign MEM[9325] = MEM[3223] + MEM[739];
assign MEM[9326] = MEM[3227] + MEM[4919];
assign MEM[9327] = MEM[3231] + MEM[6133];
assign MEM[9328] = MEM[3294] + MEM[6231];
assign MEM[9329] = MEM[3307] + MEM[5890];
assign MEM[9330] = MEM[3332] + MEM[5150];
assign MEM[9331] = MEM[3383] + MEM[4860];
assign MEM[9332] = MEM[3431] + MEM[5883];
assign MEM[9333] = MEM[3442] + MEM[5877];
assign MEM[9334] = MEM[3444] + MEM[2179];
assign MEM[9335] = MEM[3507] + MEM[5308];
assign MEM[9336] = MEM[3599] + MEM[4503];
assign MEM[9337] = MEM[3607] + MEM[5500];
assign MEM[9338] = MEM[3621] + MEM[6197];
assign MEM[9339] = MEM[3663] + MEM[4844];
assign MEM[9340] = MEM[3678] + MEM[2948];
assign MEM[9341] = MEM[3684] + MEM[6893];
assign MEM[9342] = MEM[3706] + MEM[4469];
assign MEM[9343] = MEM[3775] + MEM[5998];
assign MEM[9344] = MEM[3893] + MEM[3159];
assign MEM[9345] = MEM[3910] + MEM[3343];
assign MEM[9346] = MEM[3943] + MEM[2679];
assign MEM[9347] = MEM[3951] + MEM[4590];
assign MEM[9348] = MEM[4063] + MEM[133];
assign MEM[9349] = MEM[4102] + MEM[5293];
assign MEM[9350] = MEM[4163] + MEM[4967];
assign MEM[9351] = MEM[4166] + MEM[5981];
assign MEM[9352] = MEM[4167] + MEM[6832];
assign MEM[9353] = MEM[4213] + MEM[4772];
assign MEM[9354] = MEM[4224] + MEM[4225];
assign MEM[9355] = MEM[4302] + MEM[6054];
assign MEM[9356] = MEM[4380] + MEM[4415];
assign MEM[9357] = MEM[4406] + MEM[7038];
assign MEM[9358] = MEM[4411] + MEM[4410];
assign MEM[9359] = MEM[4426] + MEM[629];
assign MEM[9360] = MEM[4459] + MEM[5478];
assign MEM[9361] = MEM[4519] + MEM[5910];
assign MEM[9362] = MEM[4523] + MEM[1350];
assign MEM[9363] = MEM[4557] + MEM[5547];
assign MEM[9364] = MEM[4599] + MEM[2853];
assign MEM[9365] = MEM[4675] + MEM[103];
assign MEM[9366] = MEM[4730] + MEM[6126];
assign MEM[9367] = MEM[4763] + MEM[1596];
assign MEM[9368] = MEM[4781] + MEM[5866];
assign MEM[9369] = MEM[4790] + MEM[7100];
assign MEM[9370] = MEM[4806] + MEM[6951];
assign MEM[9371] = MEM[4815] + MEM[3414];
assign MEM[9372] = MEM[4845] + MEM[5599];
assign MEM[9373] = MEM[4850] + MEM[7114];
assign MEM[9374] = MEM[4911] + MEM[1837];
assign MEM[9375] = MEM[4935] + MEM[5737];
assign MEM[9376] = MEM[4942] + MEM[4429];
assign MEM[9377] = MEM[4943] + MEM[6739];
assign MEM[9378] = MEM[4998] + MEM[7054];
assign MEM[9379] = MEM[5039] + MEM[4765];
assign MEM[9380] = MEM[5108] + MEM[1110];
assign MEM[9381] = MEM[5157] + MEM[6904];
assign MEM[9382] = MEM[5186] + MEM[7134];
assign MEM[9383] = MEM[5227] + MEM[2379];
assign MEM[9384] = MEM[5229] + MEM[5397];
assign MEM[9385] = MEM[5339] + MEM[7460];
assign MEM[9386] = MEM[5406] + MEM[4029];
assign MEM[9387] = MEM[5413] + MEM[5923];
assign MEM[9388] = MEM[5583] + MEM[3759];
assign MEM[9389] = MEM[5597] + MEM[379];
assign MEM[9390] = MEM[5635] + MEM[5013];
assign MEM[9391] = MEM[5653] + MEM[4132];
assign MEM[9392] = MEM[5707] + MEM[6988];
assign MEM[9393] = MEM[5711] + MEM[2918];
assign MEM[9394] = MEM[5786] + MEM[1978];
assign MEM[9395] = MEM[5799] + MEM[5876];
assign MEM[9396] = MEM[5823] + MEM[1476];
assign MEM[9397] = MEM[5839] + MEM[1092];
assign MEM[9398] = MEM[5878] + MEM[1099];
assign MEM[9399] = MEM[5882] + MEM[942];
assign MEM[9400] = MEM[5901] + MEM[4725];
assign MEM[9401] = MEM[5942] + MEM[4882];
assign MEM[9402] = MEM[5967] + MEM[6985];
assign MEM[9403] = MEM[6015] + MEM[2099];
assign MEM[9404] = MEM[6095] + MEM[6158];
assign MEM[9405] = MEM[6118] + MEM[6953];
assign MEM[9406] = MEM[6141] + MEM[3254];
assign MEM[9407] = MEM[6165] + MEM[1251];
assign MEM[9408] = MEM[6221] + MEM[2703];
assign MEM[9409] = MEM[6239] + MEM[6995];
assign MEM[9410] = MEM[6263] + MEM[4357];
assign MEM[9411] = MEM[6692] + MEM[6915];
assign MEM[9412] = MEM[6694] + MEM[3903];
assign MEM[9413] = MEM[6779] + MEM[4878];
assign MEM[9414] = MEM[6785] + MEM[6870];
assign MEM[9415] = MEM[6797] + MEM[995];
assign MEM[9416] = MEM[6803] + MEM[7088];
assign MEM[9417] = MEM[6805] + MEM[2695];
assign MEM[9418] = MEM[6807] + MEM[7046];
assign MEM[9419] = MEM[6822] + MEM[1898];
assign MEM[9420] = MEM[6823] + MEM[7127];
assign MEM[9421] = MEM[6838] + MEM[7025];
assign MEM[9422] = MEM[6841] + MEM[7055];
assign MEM[9423] = MEM[6846] + MEM[2091];
assign MEM[9424] = MEM[6853] + MEM[6863];
assign MEM[9425] = MEM[6856] + MEM[5738];
assign MEM[9426] = MEM[6877] + MEM[6173];
assign MEM[9427] = MEM[6878] + MEM[4207];
assign MEM[9428] = MEM[6881] + MEM[7039];
assign MEM[9429] = MEM[6895] + MEM[7118];
assign MEM[9430] = MEM[6897] + MEM[6909];
assign MEM[9431] = MEM[6906] + MEM[2707];
assign MEM[9432] = MEM[6907] + MEM[7006];
assign MEM[9433] = MEM[6914] + MEM[2686];
assign MEM[9434] = MEM[6928] + MEM[6071];
assign MEM[9435] = MEM[6937] + MEM[1597];
assign MEM[9436] = MEM[6946] + MEM[3964];
assign MEM[9437] = MEM[6948] + MEM[5166];
assign MEM[9438] = MEM[6957] + MEM[7110];
assign MEM[9439] = MEM[6972] + MEM[4711];
assign MEM[9440] = MEM[6973] + MEM[6908];
assign MEM[9441] = MEM[6974] + MEM[3102];
assign MEM[9442] = MEM[6984] + MEM[6053];
assign MEM[9443] = MEM[6993] + MEM[5132];
assign MEM[9444] = MEM[7000] + MEM[7864];
assign MEM[9445] = MEM[7001] + MEM[1812];
assign MEM[9446] = MEM[7004] + MEM[3815];
assign MEM[9447] = MEM[7020] + MEM[7023];
assign MEM[9448] = MEM[7024] + MEM[3469];
assign MEM[9449] = MEM[7029] + MEM[7288];
assign MEM[9450] = MEM[7034] + MEM[7052];
assign MEM[9451] = MEM[7036] + MEM[7200];
assign MEM[9452] = MEM[7037] + MEM[7325];
assign MEM[9453] = MEM[7042] + MEM[2806];
assign MEM[9454] = MEM[7048] + MEM[1306];
assign MEM[9455] = MEM[7061] + MEM[3602];
assign MEM[9456] = MEM[7065] + MEM[7409];
assign MEM[9457] = MEM[7086] + MEM[7094];
assign MEM[9458] = MEM[7098] + MEM[7099];
assign MEM[9459] = MEM[7103] + MEM[7467];
assign MEM[9460] = MEM[7109] + MEM[7277];
assign MEM[9461] = MEM[7147] + MEM[2182];
assign MEM[9462] = MEM[7148] + MEM[7375];
assign MEM[9463] = MEM[7153] + MEM[1823];
assign MEM[9464] = MEM[7155] + MEM[7262];
assign MEM[9465] = MEM[7169] + MEM[1546];
assign MEM[9466] = MEM[7172] + MEM[7358];
assign MEM[9467] = MEM[7206] + MEM[7115];
assign MEM[9468] = MEM[7237] + MEM[7769];
assign MEM[9469] = MEM[7280] + MEM[7111];
assign MEM[9470] = MEM[7312] + MEM[4604];
assign MEM[9471] = MEM[7374] + MEM[4581];
assign MEM[9472] = MEM[7505] + MEM[3250];
assign MEM[9473] = MEM[7612] + MEM[5546];
assign MEM[9474] = MEM[7801] + MEM[5900];
assign MEM[9475] = MEM[9226] + MEM[9227];
assign MEM[9476] = MEM[23] + MEM[3149];
assign MEM[9477] = MEM[117] + MEM[5598];
assign MEM[9478] = MEM[316] + MEM[1311];
assign MEM[9479] = MEM[348] + MEM[1501];
assign MEM[9480] = MEM[350] + MEM[1706];
assign MEM[9481] = MEM[453] + MEM[511];
assign MEM[9482] = MEM[470] + MEM[7317];
assign MEM[9483] = MEM[495] + MEM[6902];
assign MEM[9484] = MEM[527] + MEM[4997];
assign MEM[9485] = MEM[532] + MEM[1930];
assign MEM[9486] = MEM[556] + MEM[2159];
assign MEM[9487] = MEM[557] + MEM[6843];
assign MEM[9488] = MEM[591] + MEM[1406];
assign MEM[9489] = MEM[603] + MEM[1430];
assign MEM[9490] = MEM[630] + MEM[1839];
assign MEM[9491] = MEM[646] + MEM[4734];
assign MEM[9492] = MEM[757] + MEM[1783];
assign MEM[9493] = MEM[957] + MEM[2954];
assign MEM[9494] = MEM[970] + MEM[4631];
assign MEM[9495] = MEM[979] + MEM[7349];
assign MEM[9496] = MEM[983] + MEM[2716];
assign MEM[9497] = MEM[1031] + MEM[1173];
assign MEM[9498] = MEM[1042] + MEM[2714];
assign MEM[9499] = MEM[1052] + MEM[3702];
assign MEM[9500] = MEM[1102] + MEM[2662];
assign MEM[9501] = MEM[1157] + MEM[1367];
assign MEM[9502] = MEM[1182] + MEM[2327];
assign MEM[9503] = MEM[1202] + MEM[3349];
assign MEM[9504] = MEM[1308] + MEM[2927];
assign MEM[9505] = MEM[1405] + MEM[1595];
assign MEM[9506] = MEM[1446] + MEM[2003];
assign MEM[9507] = MEM[1485] + MEM[6954];
assign MEM[9508] = MEM[1543] + MEM[3845];
assign MEM[9509] = MEM[1566] + MEM[2075];
assign MEM[9510] = MEM[1612] + MEM[5299];
assign MEM[9511] = MEM[1643] + MEM[7106];
assign MEM[9512] = MEM[1644] + MEM[4110];
assign MEM[9513] = MEM[1682] + MEM[8131];
assign MEM[9514] = MEM[1821] + MEM[3447];
assign MEM[9515] = MEM[1886] + MEM[830];
assign MEM[9516] = MEM[1887] + MEM[4917];
assign MEM[9517] = MEM[1901] + MEM[2706];
assign MEM[9518] = MEM[1938] + MEM[1939];
assign MEM[9519] = MEM[2005] + MEM[6976];
assign MEM[9520] = MEM[2059] + MEM[2422];
assign MEM[9521] = MEM[2063] + MEM[5187];
assign MEM[9522] = MEM[2147] + MEM[3295];
assign MEM[9523] = MEM[2172] + MEM[7371];
assign MEM[9524] = MEM[2231] + MEM[3059];
assign MEM[9525] = MEM[2255] + MEM[4565];
assign MEM[9526] = MEM[2351] + MEM[5135];
assign MEM[9527] = MEM[2455] + MEM[5286];
assign MEM[9528] = MEM[2645] + MEM[6968];
assign MEM[9529] = MEM[2755] + MEM[4814];
assign MEM[9530] = MEM[2779] + MEM[6246];
assign MEM[9531] = MEM[2879] + MEM[3078];
assign MEM[9532] = MEM[2902] + MEM[4852];
assign MEM[9533] = MEM[2932] + MEM[6922];
assign MEM[9534] = MEM[2981] + MEM[6913];
assign MEM[9535] = MEM[2994] + MEM[5261];
assign MEM[9536] = MEM[3036] + MEM[671];
assign MEM[9537] = MEM[3068] + MEM[5445];
assign MEM[9538] = MEM[3086] + MEM[7074];
assign MEM[9539] = MEM[3101] + MEM[1307];
assign MEM[9540] = MEM[3156] + MEM[6923];
assign MEM[9541] = MEM[3166] + MEM[5028];
assign MEM[9542] = MEM[3188] + MEM[4910];
assign MEM[9543] = MEM[3197] + MEM[5276];
assign MEM[9544] = MEM[3236] + MEM[5515];
assign MEM[9545] = MEM[3381] + MEM[5709];
assign MEM[9546] = MEM[3411] + MEM[7075];
assign MEM[9547] = MEM[3426] + MEM[3434];
assign MEM[9548] = MEM[3468] + MEM[7179];
assign MEM[9549] = MEM[3722] + MEM[7254];
assign MEM[9550] = MEM[3786] + MEM[3326];
assign MEM[9551] = MEM[3787] + MEM[5639];
assign MEM[9552] = MEM[3855] + MEM[4013];
assign MEM[9553] = MEM[3859] + MEM[7122];
assign MEM[9554] = MEM[3898] + MEM[2572];
assign MEM[9555] = MEM[3916] + MEM[5007];
assign MEM[9556] = MEM[3933] + MEM[5221];
assign MEM[9557] = MEM[3957] + MEM[1285];
assign MEM[9558] = MEM[4012] + MEM[7062];
assign MEM[9559] = MEM[4068] + MEM[7159];
assign MEM[9560] = MEM[4109] + MEM[1690];
assign MEM[9561] = MEM[4118] + MEM[1996];
assign MEM[9562] = MEM[4151] + MEM[4190];
assign MEM[9563] = MEM[4174] + MEM[5775];
assign MEM[9564] = MEM[4187] + MEM[7084];
assign MEM[9565] = MEM[4210] + MEM[7763];
assign MEM[9566] = MEM[4236] + MEM[4686];
assign MEM[9567] = MEM[4438] + MEM[7119];
assign MEM[9568] = MEM[4442] + MEM[5459];
assign MEM[9569] = MEM[4479] + MEM[2295];
assign MEM[9570] = MEM[4506] + MEM[788];
assign MEM[9571] = MEM[4571] + MEM[7059];
assign MEM[9572] = MEM[4613] + MEM[6876];
assign MEM[9573] = MEM[4627] + MEM[5644];
assign MEM[9574] = MEM[4685] + MEM[1199];
assign MEM[9575] = MEM[4779] + MEM[4069];
assign MEM[9576] = MEM[4794] + MEM[7051];
assign MEM[9577] = MEM[4829] + MEM[1204];
assign MEM[9578] = MEM[4894] + MEM[4903];
assign MEM[9579] = MEM[4991] + MEM[7281];
assign MEM[9580] = MEM[4999] + MEM[5301];
assign MEM[9581] = MEM[5030] + MEM[5095];
assign MEM[9582] = MEM[5071] + MEM[2989];
assign MEM[9583] = MEM[5127] + MEM[3047];
assign MEM[9584] = MEM[5215] + MEM[7138];
assign MEM[9585] = MEM[5278] + MEM[6774];
assign MEM[9586] = MEM[5395] + MEM[5853];
assign MEM[9587] = MEM[5450] + MEM[3300];
assign MEM[9588] = MEM[5535] + MEM[6938];
assign MEM[9589] = MEM[5591] + MEM[2238];
assign MEM[9590] = MEM[5690] + MEM[5791];
assign MEM[9591] = MEM[5746] + MEM[1293];
assign MEM[9592] = MEM[5759] + MEM[7139];
assign MEM[9593] = MEM[5796] + MEM[3007];
assign MEM[9594] = MEM[5907] + MEM[5313];
assign MEM[9595] = MEM[5922] + MEM[7083];
assign MEM[9596] = MEM[5932] + MEM[7072];
assign MEM[9597] = MEM[5963] + MEM[2612];
assign MEM[9598] = MEM[6102] + MEM[6980];
assign MEM[9599] = MEM[6109] + MEM[3375];
assign MEM[9600] = MEM[6163] + MEM[7027];
assign MEM[9601] = MEM[6166] + MEM[1036];
assign MEM[9602] = MEM[6254] + MEM[4083];
assign MEM[9603] = MEM[6262] + MEM[5757];
assign MEM[9604] = MEM[6806] + MEM[710];
assign MEM[9605] = MEM[6810] + MEM[6930];
assign MEM[9606] = MEM[6901] + MEM[5647];
assign MEM[9607] = MEM[6949] + MEM[325];
assign MEM[9608] = MEM[6959] + MEM[2227];
assign MEM[9609] = MEM[6964] + MEM[1279];
assign MEM[9610] = MEM[6966] + MEM[1541];
assign MEM[9611] = MEM[6969] + MEM[2098];
assign MEM[9612] = MEM[6996] + MEM[835];
assign MEM[9613] = MEM[6998] + MEM[3421];
assign MEM[9614] = MEM[6999] + MEM[5550];
assign MEM[9615] = MEM[7003] + MEM[2660];
assign MEM[9616] = MEM[7011] + MEM[5774];
assign MEM[9617] = MEM[7013] + MEM[7104];
assign MEM[9618] = MEM[7019] + MEM[7786];
assign MEM[9619] = MEM[7028] + MEM[7201];
assign MEM[9620] = MEM[7031] + MEM[612];
assign MEM[9621] = MEM[7032] + MEM[1634];
assign MEM[9622] = MEM[7043] + MEM[2036];
assign MEM[9623] = MEM[7053] + MEM[4789];
assign MEM[9624] = MEM[7057] + MEM[2565];
assign MEM[9625] = MEM[7060] + MEM[4134];
assign MEM[9626] = MEM[7076] + MEM[7345];
assign MEM[9627] = MEM[7096] + MEM[7357];
assign MEM[9628] = MEM[7097] + MEM[4514];
assign MEM[9629] = MEM[7105] + MEM[2093];
assign MEM[9630] = MEM[7120] + MEM[7197];
assign MEM[9631] = MEM[7121] + MEM[14];
assign MEM[9632] = MEM[7144] + MEM[2122];
assign MEM[9633] = MEM[7149] + MEM[5181];
assign MEM[9634] = MEM[7152] + MEM[7389];
assign MEM[9635] = MEM[7161] + MEM[5925];
assign MEM[9636] = MEM[7167] + MEM[3661];
assign MEM[9637] = MEM[7171] + MEM[4283];
assign MEM[9638] = MEM[7173] + MEM[7707];
assign MEM[9639] = MEM[7175] + MEM[2789];
assign MEM[9640] = MEM[7176] + MEM[7339];
assign MEM[9641] = MEM[7177] + MEM[7578];
assign MEM[9642] = MEM[7180] + MEM[628];
assign MEM[9643] = MEM[7199] + MEM[963];
assign MEM[9644] = MEM[7204] + MEM[7116];
assign MEM[9645] = MEM[7212] + MEM[5003];
assign MEM[9646] = MEM[7213] + MEM[7323];
assign MEM[9647] = MEM[7219] + MEM[7191];
assign MEM[9648] = MEM[7238] + MEM[2995];
assign MEM[9649] = MEM[7273] + MEM[8084];
assign MEM[9650] = MEM[7334] + MEM[7817];
assign MEM[9651] = MEM[7352] + MEM[7860];
assign MEM[9652] = MEM[7366] + MEM[1749];
assign MEM[9653] = MEM[7373] + MEM[6924];
assign MEM[9654] = MEM[7376] + MEM[7600];
assign MEM[9655] = MEM[7381] + MEM[6801];
assign MEM[9656] = MEM[7421] + MEM[741];
assign MEM[9657] = MEM[7531] + MEM[7151];
assign MEM[9658] = MEM[7536] + MEM[7560];
assign MEM[9659] = MEM[7566] + MEM[4892];
assign MEM[9660] = MEM[7841] + MEM[4427];
assign MEM[9661] = MEM[7856] + MEM[6107];
assign MEM[9662] = MEM[7865] + MEM[7422];
assign MEM[9663] = MEM[7872] + MEM[8048];
assign MEM[9664] = MEM[8028] + MEM[8134];
assign MEM[9665] = MEM[8132] + MEM[791];
assign MEM[9666] = MEM[222] + MEM[5285];
assign MEM[9667] = MEM[223] + MEM[588];
assign MEM[9668] = MEM[284] + MEM[311];
assign MEM[9669] = MEM[294] + MEM[5235];
assign MEM[9670] = MEM[371] + MEM[5094];
assign MEM[9671] = MEM[455] + MEM[6967];
assign MEM[9672] = MEM[548] + MEM[4926];
assign MEM[9673] = MEM[567] + MEM[4842];
assign MEM[9674] = MEM[570] + MEM[3807];
assign MEM[9675] = MEM[744] + MEM[7771];
assign MEM[9676] = MEM[748] + MEM[2637];
assign MEM[9677] = MEM[778] + MEM[5054];
assign MEM[9678] = MEM[781] + MEM[7278];
assign MEM[9679] = MEM[819] + MEM[2070];
assign MEM[9680] = MEM[956] + MEM[1716];
assign MEM[9681] = MEM[974] + MEM[2202];
assign MEM[9682] = MEM[1020] + MEM[7315];
assign MEM[9683] = MEM[1091] + MEM[5143];
assign MEM[9684] = MEM[1150] + MEM[1578];
assign MEM[9685] = MEM[1162] + MEM[4621];
assign MEM[9686] = MEM[1180] + MEM[5645];
assign MEM[9687] = MEM[1214] + MEM[5589];
assign MEM[9688] = MEM[1268] + MEM[2294];
assign MEM[9689] = MEM[1286] + MEM[5444];
assign MEM[9690] = MEM[1310] + MEM[5782];
assign MEM[9691] = MEM[1325] + MEM[3532];
assign MEM[9692] = MEM[1527] + MEM[2427];
assign MEM[9693] = MEM[1530] + MEM[5574];
assign MEM[9694] = MEM[1539] + MEM[1855];
assign MEM[9695] = MEM[1579] + MEM[7328];
assign MEM[9696] = MEM[1607] + MEM[2602];
assign MEM[9697] = MEM[1653] + MEM[2687];
assign MEM[9698] = MEM[1654] + MEM[5988];
assign MEM[9699] = MEM[1668] + MEM[7320];
assign MEM[9700] = MEM[1679] + MEM[5830];
assign MEM[9701] = MEM[1733] + MEM[5485];
assign MEM[9702] = MEM[1815] + MEM[7257];
assign MEM[9703] = MEM[1883] + MEM[7090];
assign MEM[9704] = MEM[1884] + MEM[1395];
assign MEM[9705] = MEM[1899] + MEM[7026];
assign MEM[9706] = MEM[1914] + MEM[5542];
assign MEM[9707] = MEM[1965] + MEM[3643];
assign MEM[9708] = MEM[1971] + MEM[2470];
assign MEM[9709] = MEM[1988] + MEM[3541];
assign MEM[9710] = MEM[2054] + MEM[3220];
assign MEM[9711] = MEM[2203] + MEM[2692];
assign MEM[9712] = MEM[2212] + MEM[7326];
assign MEM[9713] = MEM[2271] + MEM[2650];
assign MEM[9714] = MEM[2276] + MEM[4186];
assign MEM[9715] = MEM[2278] + MEM[3242];
assign MEM[9716] = MEM[2370] + MEM[7695];
assign MEM[9717] = MEM[2373] + MEM[6135];
assign MEM[9718] = MEM[2402] + MEM[7395];
assign MEM[9719] = MEM[2420] + MEM[3158];
assign MEM[9720] = MEM[2615] + MEM[2807];
assign MEM[9721] = MEM[2701] + MEM[5067];
assign MEM[9722] = MEM[2715] + MEM[2606];
assign MEM[9723] = MEM[2734] + MEM[5123];
assign MEM[9724] = MEM[2767] + MEM[4693];
assign MEM[9725] = MEM[2795] + MEM[3494];
assign MEM[9726] = MEM[2971] + MEM[2733];
assign MEM[9727] = MEM[3082] + MEM[5543];
assign MEM[9728] = MEM[3087] + MEM[7252];
assign MEM[9729] = MEM[3126] + MEM[3719];
assign MEM[9730] = MEM[3270] + MEM[4111];
assign MEM[9731] = MEM[3301] + MEM[2583];
assign MEM[9732] = MEM[3390] + MEM[7523];
assign MEM[9733] = MEM[3485] + MEM[4407];
assign MEM[9734] = MEM[3517] + MEM[3835];
assign MEM[9735] = MEM[3639] + MEM[7216];
assign MEM[9736] = MEM[3677] + MEM[4294];
assign MEM[9737] = MEM[3695] + MEM[485];
assign MEM[9738] = MEM[3747] + MEM[7091];
assign MEM[9739] = MEM[3762] + MEM[5911];
assign MEM[9740] = MEM[3907] + MEM[5312];
assign MEM[9741] = MEM[3940] + MEM[3948];
assign MEM[9742] = MEM[4044] + MEM[7140];
assign MEM[9743] = MEM[4046] + MEM[7651];
assign MEM[9744] = MEM[4126] + MEM[5165];
assign MEM[9745] = MEM[4178] + MEM[7354];
assign MEM[9746] = MEM[4191] + MEM[3348];
assign MEM[9747] = MEM[4205] + MEM[7300];
assign MEM[9748] = MEM[4262] + MEM[5219];
assign MEM[9749] = MEM[4292] + MEM[5715];
assign MEM[9750] = MEM[4303] + MEM[7063];
assign MEM[9751] = MEM[4309] + MEM[7306];
assign MEM[9752] = MEM[4342] + MEM[4787];
assign MEM[9753] = MEM[4367] + MEM[5771];
assign MEM[9754] = MEM[4412] + MEM[2127];
assign MEM[9755] = MEM[4435] + MEM[5426];
assign MEM[9756] = MEM[4532] + MEM[6178];
assign MEM[9757] = MEM[4546] + MEM[4547];
assign MEM[9758] = MEM[4559] + MEM[7321];
assign MEM[9759] = MEM[4589] + MEM[7335];
assign MEM[9760] = MEM[4638] + MEM[4995];
assign MEM[9761] = MEM[4666] + MEM[7142];
assign MEM[9762] = MEM[4731] + MEM[3395];
assign MEM[9763] = MEM[4821] + MEM[3598];
assign MEM[9764] = MEM[4828] + MEM[5498];
assign MEM[9765] = MEM[4839] + MEM[7605];
assign MEM[9766] = MEM[4854] + MEM[5666];
assign MEM[9767] = MEM[4895] + MEM[6983];
assign MEM[9768] = MEM[4954] + MEM[3461];
assign MEM[9769] = MEM[4956] + MEM[367];
assign MEM[9770] = MEM[5151] + MEM[4963];
assign MEM[9771] = MEM[5182] + MEM[6181];
assign MEM[9772] = MEM[5199] + MEM[7272];
assign MEM[9773] = MEM[5203] + MEM[5642];
assign MEM[9774] = MEM[5220] + MEM[7245];
assign MEM[9775] = MEM[5234] + MEM[1149];
assign MEM[9776] = MEM[5267] + MEM[7420];
assign MEM[9777] = MEM[5314] + MEM[6078];
assign MEM[9778] = MEM[5374] + MEM[6975];
assign MEM[9779] = MEM[5381] + MEM[2541];
assign MEM[9780] = MEM[5454] + MEM[7283];
assign MEM[9781] = MEM[5467] + MEM[7126];
assign MEM[9782] = MEM[5501] + MEM[7108];
assign MEM[9783] = MEM[5503] + MEM[7209];
assign MEM[9784] = MEM[5517] + MEM[6230];
assign MEM[9785] = MEM[5522] + MEM[5548];
assign MEM[9786] = MEM[5523] + MEM[5534];
assign MEM[9787] = MEM[5563] + MEM[7146];
assign MEM[9788] = MEM[5565] + MEM[7211];
assign MEM[9789] = MEM[5566] + MEM[1332];
assign MEM[9790] = MEM[5579] + MEM[7385];
assign MEM[9791] = MEM[5714] + MEM[1319];
assign MEM[9792] = MEM[5730] + MEM[7298];
assign MEM[9793] = MEM[5924] + MEM[7507];
assign MEM[9794] = MEM[5958] + MEM[7217];
assign MEM[9795] = MEM[5978] + MEM[869];
assign MEM[9796] = MEM[6047] + MEM[6945];
assign MEM[9797] = MEM[6111] + MEM[2157];
assign MEM[9798] = MEM[6134] + MEM[6174];
assign MEM[9799] = MEM[6180] + MEM[7318];
assign MEM[9800] = MEM[6189] + MEM[3175];
assign MEM[9801] = MEM[6270] + MEM[7214];
assign MEM[9802] = MEM[7047] + MEM[7137];
assign MEM[9803] = MEM[7073] + MEM[3043];
assign MEM[9804] = MEM[7087] + MEM[7486];
assign MEM[9805] = MEM[7095] + MEM[7247];
assign MEM[9806] = MEM[7101] + MEM[595];
assign MEM[9807] = MEM[7102] + MEM[7471];
assign MEM[9808] = MEM[7107] + MEM[5667];
assign MEM[9809] = MEM[7112] + MEM[7482];
assign MEM[9810] = MEM[7123] + MEM[7310];
assign MEM[9811] = MEM[7124] + MEM[7224];
assign MEM[9812] = MEM[7129] + MEM[7499];
assign MEM[9813] = MEM[7130] + MEM[5451];
assign MEM[9814] = MEM[7133] + MEM[562];
assign MEM[9815] = MEM[7154] + MEM[7311];
assign MEM[9816] = MEM[7162] + MEM[7364];
assign MEM[9817] = MEM[7205] + MEM[5682];
assign MEM[9818] = MEM[7208] + MEM[5997];
assign MEM[9819] = MEM[7210] + MEM[7276];
assign MEM[9820] = MEM[7218] + MEM[5342];
assign MEM[9821] = MEM[7236] + MEM[5270];
assign MEM[9822] = MEM[7241] + MEM[7];
assign MEM[9823] = MEM[7242] + MEM[4580];
assign MEM[9824] = MEM[7246] + MEM[4402];
assign MEM[9825] = MEM[7261] + MEM[7481];
assign MEM[9826] = MEM[7268] + MEM[3218];
assign MEM[9827] = MEM[7269] + MEM[5541];
assign MEM[9828] = MEM[7271] + MEM[7340];
assign MEM[9829] = MEM[7285] + MEM[7304];
assign MEM[9830] = MEM[7287] + MEM[7510];
assign MEM[9831] = MEM[7293] + MEM[5189];
assign MEM[9832] = MEM[7297] + MEM[4986];
assign MEM[9833] = MEM[7301] + MEM[501];
assign MEM[9834] = MEM[7302] + MEM[4290];
assign MEM[9835] = MEM[7314] + MEM[7327];
assign MEM[9836] = MEM[7322] + MEM[5806];
assign MEM[9837] = MEM[7332] + MEM[7244];
assign MEM[9838] = MEM[7338] + MEM[7392];
assign MEM[9839] = MEM[7351] + MEM[7166];
assign MEM[9840] = MEM[7355] + MEM[7545];
assign MEM[9841] = MEM[7367] + MEM[7541];
assign MEM[9842] = MEM[7369] + MEM[4052];
assign MEM[9843] = MEM[7372] + MEM[7520];
assign MEM[9844] = MEM[7383] + MEM[7432];
assign MEM[9845] = MEM[7384] + MEM[2469];
assign MEM[9846] = MEM[7413] + MEM[2222];
assign MEM[9847] = MEM[7428] + MEM[7739];
assign MEM[9848] = MEM[7429] + MEM[7589];
assign MEM[9849] = MEM[7435] + MEM[4014];
assign MEM[9850] = MEM[7443] + MEM[7472];
assign MEM[9851] = MEM[7451] + MEM[7690];
assign MEM[9852] = MEM[7470] + MEM[7457];
assign MEM[9853] = MEM[7491] + MEM[5173];
assign MEM[9854] = MEM[7495] + MEM[7480];
assign MEM[9855] = MEM[7508] + MEM[7625];
assign MEM[9856] = MEM[7530] + MEM[7743];
assign MEM[9857] = MEM[7539] + MEM[1882];
assign MEM[9858] = MEM[7643] + MEM[7407];
assign MEM[9859] = MEM[7697] + MEM[7775];
assign MEM[9860] = MEM[7797] + MEM[4084];
assign MEM[9861] = MEM[7808] + MEM[7883];
assign MEM[9862] = MEM[7843] + MEM[7842];
assign MEM[9863] = MEM[7958] + MEM[7497];
assign MEM[9864] = MEM[8467] + MEM[7552];
assign MEM[9865] = MEM[9857] + MEM[7706];
assign MEM[9866] = MEM[9861] + MEM[5042];
assign MEM[9867] = MEM[69] + MEM[5325];
assign MEM[9868] = MEM[317] + MEM[3851];
assign MEM[9869] = MEM[483] + MEM[3306];
assign MEM[9870] = MEM[598] + MEM[1010];
assign MEM[9871] = MEM[627] + MEM[8337];
assign MEM[9872] = MEM[727] + MEM[1318];
assign MEM[9873] = MEM[853] + MEM[1747];
assign MEM[9874] = MEM[911] + MEM[1660];
assign MEM[9875] = MEM[975] + MEM[2812];
assign MEM[9876] = MEM[991] + MEM[2387];
assign MEM[9877] = MEM[1053] + MEM[5303];
assign MEM[9878] = MEM[1061] + MEM[4282];
assign MEM[9879] = MEM[1098] + MEM[7386];
assign MEM[9880] = MEM[1111] + MEM[1002];
assign MEM[9881] = MEM[1218] + MEM[7540];
assign MEM[9882] = MEM[1404] + MEM[7243];
assign MEM[9883] = MEM[1468] + MEM[1724];
assign MEM[9884] = MEM[1474] + MEM[7461];
assign MEM[9885] = MEM[1482] + MEM[4876];
assign MEM[9886] = MEM[1581] + MEM[5422];
assign MEM[9887] = MEM[1615] + MEM[1255];
assign MEM[9888] = MEM[1629] + MEM[7439];
assign MEM[9889] = MEM[1732] + MEM[7390];
assign MEM[9890] = MEM[1955] + MEM[4351];
assign MEM[9891] = MEM[2102] + MEM[4541];
assign MEM[9892] = MEM[2162] + MEM[2386];
assign MEM[9893] = MEM[2163] + MEM[7291];
assign MEM[9894] = MEM[2170] + MEM[2171];
assign MEM[9895] = MEM[2178] + MEM[3463];
assign MEM[9896] = MEM[2194] + MEM[3404];
assign MEM[9897] = MEM[2259] + MEM[2967];
assign MEM[9898] = MEM[2275] + MEM[1669];
assign MEM[9899] = MEM[2341] + MEM[7689];
assign MEM[9900] = MEM[2423] + MEM[2850];
assign MEM[9901] = MEM[2595] + MEM[986];
assign MEM[9902] = MEM[2626] + MEM[7248];
assign MEM[9903] = MEM[2655] + MEM[7353];
assign MEM[9904] = MEM[2773] + MEM[5133];
assign MEM[9905] = MEM[2781] + MEM[7240];
assign MEM[9906] = MEM[2787] + MEM[2794];
assign MEM[9907] = MEM[2852] + MEM[5050];
assign MEM[9908] = MEM[2926] + MEM[7549];
assign MEM[9909] = MEM[3023] + MEM[3027];
assign MEM[9910] = MEM[3061] + MEM[4983];
assign MEM[9911] = MEM[3083] + MEM[7368];
assign MEM[9912] = MEM[3141] + MEM[4587];
assign MEM[9913] = MEM[3221] + MEM[5447];
assign MEM[9914] = MEM[3237] + MEM[599];
assign MEM[9915] = MEM[3283] + MEM[4972];
assign MEM[9916] = MEM[3410] + MEM[407];
assign MEM[9917] = MEM[3429] + MEM[7745];
assign MEM[9918] = MEM[3467] + MEM[5346];
assign MEM[9919] = MEM[3535] + MEM[5069];
assign MEM[9920] = MEM[3570] + MEM[6255];
assign MEM[9921] = MEM[3662] + MEM[4682];
assign MEM[9922] = MEM[3703] + MEM[7574];
assign MEM[9923] = MEM[3788] + MEM[7537];
assign MEM[9924] = MEM[3838] + MEM[7292];
assign MEM[9925] = MEM[3860] + MEM[7377];
assign MEM[9926] = MEM[4005] + MEM[4902];
assign MEM[9927] = MEM[4183] + MEM[4420];
assign MEM[9928] = MEM[4263] + MEM[5740];
assign MEM[9929] = MEM[4275] + MEM[6070];
assign MEM[9930] = MEM[4323] + MEM[7622];
assign MEM[9931] = MEM[4356] + MEM[7330];
assign MEM[9932] = MEM[4476] + MEM[7483];
assign MEM[9933] = MEM[4478] + MEM[4890];
assign MEM[9934] = MEM[4578] + MEM[4331];
assign MEM[9935] = MEM[4654] + MEM[7380];
assign MEM[9936] = MEM[4660] + MEM[6030];
assign MEM[9937] = MEM[4710] + MEM[3196];
assign MEM[9938] = MEM[4724] + MEM[5210];
assign MEM[9939] = MEM[4733] + MEM[5326];
assign MEM[9940] = MEM[4855] + MEM[5412];
assign MEM[9941] = MEM[4868] + MEM[7391];
assign MEM[9942] = MEM[4877] + MEM[4989];
assign MEM[9943] = MEM[5011] + MEM[7145];
assign MEM[9944] = MEM[5019] + MEM[4362];
assign MEM[9945] = MEM[5035] + MEM[7496];
assign MEM[9946] = MEM[5218] + MEM[5637];
assign MEM[9947] = MEM[5239] + MEM[7308];
assign MEM[9948] = MEM[5343] + MEM[7414];
assign MEM[9949] = MEM[5458] + MEM[7430];
assign MEM[9950] = MEM[5492] + MEM[2646];
assign MEM[9951] = MEM[5516] + MEM[7597];
assign MEM[9952] = MEM[5580] + MEM[7419];
assign MEM[9953] = MEM[5659] + MEM[3333];
assign MEM[9954] = MEM[5684] + MEM[1555];
assign MEM[9955] = MEM[5698] + MEM[7365];
assign MEM[9956] = MEM[5748] + MEM[7324];
assign MEM[9957] = MEM[5751] + MEM[8177];
assign MEM[9958] = MEM[5855] + MEM[1646];
assign MEM[9959] = MEM[5972] + MEM[7664];
assign MEM[9960] = MEM[6110] + MEM[7616];
assign MEM[9961] = MEM[6142] + MEM[7239];
assign MEM[9962] = MEM[6182] + MEM[7785];
assign MEM[9963] = MEM[7143] + MEM[4637];
assign MEM[9964] = MEM[7178] + MEM[7794];
assign MEM[9965] = MEM[7198] + MEM[7548];
assign MEM[9966] = MEM[7207] + MEM[7393];
assign MEM[9967] = MEM[7215] + MEM[2531];
assign MEM[9968] = MEM[7234] + MEM[7294];
assign MEM[9969] = MEM[7235] + MEM[7813];
assign MEM[9970] = MEM[7249] + MEM[8029];
assign MEM[9971] = MEM[7256] + MEM[7289];
assign MEM[9972] = MEM[7270] + MEM[1170];
assign MEM[9973] = MEM[7275] + MEM[7511];
assign MEM[9974] = MEM[7282] + MEM[7378];
assign MEM[9975] = MEM[7299] + MEM[7316];
assign MEM[9976] = MEM[7305] + MEM[7598];
assign MEM[9977] = MEM[7307] + MEM[4719];
assign MEM[9978] = MEM[7337] + MEM[582];
assign MEM[9979] = MEM[7343] + MEM[998];
assign MEM[9980] = MEM[7344] + MEM[7454];
assign MEM[9981] = MEM[7350] + MEM[7479];
assign MEM[9982] = MEM[7359] + MEM[2103];
assign MEM[9983] = MEM[7370] + MEM[7538];
assign MEM[9984] = MEM[7382] + MEM[7661];
assign MEM[9985] = MEM[7387] + MEM[7403];
assign MEM[9986] = MEM[7388] + MEM[7614];
assign MEM[9987] = MEM[7394] + MEM[1013];
assign MEM[9988] = MEM[7410] + MEM[1611];
assign MEM[9989] = MEM[7423] + MEM[3939];
assign MEM[9990] = MEM[7424] + MEM[4148];
assign MEM[9991] = MEM[7431] + MEM[1050];
assign MEM[9992] = MEM[7434] + MEM[8107];
assign MEM[9993] = MEM[7438] + MEM[4539];
assign MEM[9994] = MEM[7441] + MEM[7478];
assign MEM[9995] = MEM[7442] + MEM[7455];
assign MEM[9996] = MEM[7452] + MEM[7512];
assign MEM[9997] = MEM[7462] + MEM[7572];
assign MEM[9998] = MEM[7468] + MEM[7727];
assign MEM[9999] = MEM[7469] + MEM[2067];
assign MEM[10000] = MEM[7476] + MEM[5407];
assign MEM[10001] = MEM[7477] + MEM[7704];
assign MEM[10002] = MEM[7489] + MEM[7604];
assign MEM[10003] = MEM[7502] + MEM[7744];
assign MEM[10004] = MEM[7503] + MEM[7965];
assign MEM[10005] = MEM[7518] + MEM[7595];
assign MEM[10006] = MEM[7524] + MEM[191];
assign MEM[10007] = MEM[7528] + MEM[7723];
assign MEM[10008] = MEM[7534] + MEM[7547];
assign MEM[10009] = MEM[7546] + MEM[8005];
assign MEM[10010] = MEM[7550] + MEM[7593];
assign MEM[10011] = MEM[7551] + MEM[7573];
assign MEM[10012] = MEM[7562] + MEM[7620];
assign MEM[10013] = MEM[7567] + MEM[7618];
assign MEM[10014] = MEM[7570] + MEM[7571];
assign MEM[10015] = MEM[7576] + MEM[8283];
assign MEM[10016] = MEM[7594] + MEM[7225];
assign MEM[10017] = MEM[7599] + MEM[7787];
assign MEM[10018] = MEM[7601] + MEM[7862];
assign MEM[10019] = MEM[7603] + MEM[7610];
assign MEM[10020] = MEM[7606] + MEM[3107];
assign MEM[10021] = MEM[7607] + MEM[8026];
assign MEM[10022] = MEM[7609] + MEM[7615];
assign MEM[10023] = MEM[7611] + MEM[7944];
assign MEM[10024] = MEM[7621] + MEM[7613];
assign MEM[10025] = MEM[7623] + MEM[8100];
assign MEM[10026] = MEM[7633] + MEM[7852];
assign MEM[10027] = MEM[7645] + MEM[5790];
assign MEM[10028] = MEM[7646] + MEM[2860];
assign MEM[10029] = MEM[7657] + MEM[8184];
assign MEM[10030] = MEM[7668] + MEM[8191];
assign MEM[10031] = MEM[7676] + MEM[493];
assign MEM[10032] = MEM[7684] + MEM[8049];
assign MEM[10033] = MEM[7701] + MEM[8413];
assign MEM[10034] = MEM[7715] + MEM[8493];
assign MEM[10035] = MEM[7731] + MEM[7768];
assign MEM[10036] = MEM[7733] + MEM[7962];
assign MEM[10037] = MEM[7746] + MEM[7945];
assign MEM[10038] = MEM[7756] + MEM[4279];
assign MEM[10039] = MEM[7757] + MEM[7737];
assign MEM[10040] = MEM[7760] + MEM[8033];
assign MEM[10041] = MEM[7782] + MEM[8066];
assign MEM[10042] = MEM[7789] + MEM[7790];
assign MEM[10043] = MEM[7800] + MEM[7824];
assign MEM[10044] = MEM[7827] + MEM[7501];
assign MEM[10045] = MEM[7836] + MEM[2298];
assign MEM[10046] = MEM[7837] + MEM[7631];
assign MEM[10047] = MEM[7839] + MEM[2047];
assign MEM[10048] = MEM[7854] + MEM[7592];
assign MEM[10049] = MEM[7882] + MEM[2154];
assign MEM[10050] = MEM[7916] + MEM[7295];
assign MEM[10051] = MEM[7963] + MEM[868];
assign MEM[10052] = MEM[7976] + MEM[8116];
assign MEM[10053] = MEM[7998] + MEM[7869];
assign MEM[10054] = MEM[8045] + MEM[7735];
assign MEM[10055] = MEM[8055] + MEM[5236];
assign MEM[10056] = MEM[8108] + MEM[8218];
assign MEM[10057] = MEM[8109] + MEM[7692];
assign MEM[10058] = MEM[8112] + MEM[7711];
assign MEM[10059] = MEM[8133] + MEM[7602];
assign MEM[10060] = MEM[8650] + MEM[596];
assign MEM[10061] = MEM[9907] + MEM[7561];
assign MEM[10062] = MEM[516] + MEM[4123];
assign MEM[10063] = MEM[586] + MEM[7654];
assign MEM[10064] = MEM[623] + MEM[7628];
assign MEM[10065] = MEM[745] + MEM[4455];
assign MEM[10066] = MEM[831] + MEM[2207];
assign MEM[10067] = MEM[860] + MEM[1277];
assign MEM[10068] = MEM[966] + MEM[7747];
assign MEM[10069] = MEM[993] + MEM[992];
assign MEM[10070] = MEM[1302] + MEM[8148];
assign MEM[10071] = MEM[1359] + MEM[7847];
assign MEM[10072] = MEM[1411] + MEM[7975];
assign MEM[10073] = MEM[1435] + MEM[7791];
assign MEM[10074] = MEM[1470] + MEM[5700];
assign MEM[10075] = MEM[1598] + MEM[3252];
assign MEM[10076] = MEM[1635] + MEM[2875];
assign MEM[10077] = MEM[1692] + MEM[7464];
assign MEM[10078] = MEM[1710] + MEM[726];
assign MEM[10079] = MEM[1742] + MEM[5692];
assign MEM[10080] = MEM[1798] + MEM[7627];
assign MEM[10081] = MEM[1845] + MEM[3924];
assign MEM[10082] = MEM[1918] + MEM[647];
assign MEM[10083] = MEM[2012] + MEM[7519];
assign MEM[10084] = MEM[2074] + MEM[5995];
assign MEM[10085] = MEM[2082] + MEM[7458];
assign MEM[10086] = MEM[2158] + MEM[1589];
assign MEM[10087] = MEM[2254] + MEM[8053];
assign MEM[10088] = MEM[2286] + MEM[7881];
assign MEM[10089] = MEM[2468] + MEM[7885];
assign MEM[10090] = MEM[2511] + MEM[7970];
assign MEM[10091] = MEM[2658] + MEM[7720];
assign MEM[10092] = MEM[2790] + MEM[7517];
assign MEM[10093] = MEM[2847] + MEM[2815];
assign MEM[10094] = MEM[2861] + MEM[7725];
assign MEM[10095] = MEM[3031] + MEM[7698];
assign MEM[10096] = MEM[3042] + MEM[7796];
assign MEM[10097] = MEM[3286] + MEM[7919];
assign MEM[10098] = MEM[3509] + MEM[7802];
assign MEM[10099] = MEM[3556] + MEM[7580];
assign MEM[10100] = MEM[3572] + MEM[5214];
assign MEM[10101] = MEM[3690] + MEM[4237];
assign MEM[10102] = MEM[3725] + MEM[7678];
assign MEM[10103] = MEM[3749] + MEM[7868];
assign MEM[10104] = MEM[3794] + MEM[4031];
assign MEM[10105] = MEM[3806] + MEM[7703];
assign MEM[10106] = MEM[3823] + MEM[8169];
assign MEM[10107] = MEM[3834] + MEM[8036];
assign MEM[10108] = MEM[3935] + MEM[7988];
assign MEM[10109] = MEM[3975] + MEM[7649];
assign MEM[10110] = MEM[4060] + MEM[4359];
assign MEM[10111] = MEM[4139] + MEM[7329];
assign MEM[10112] = MEM[4182] + MEM[7873];
assign MEM[10113] = MEM[4222] + MEM[8098];
assign MEM[10114] = MEM[4365] + MEM[4510];
assign MEM[10115] = MEM[4447] + MEM[4540];
assign MEM[10116] = MEM[4467] + MEM[7279];
assign MEM[10117] = MEM[4472] + MEM[4473];
assign MEM[10118] = MEM[4474] + MEM[10117];
assign MEM[10119] = MEM[4477] + MEM[4538];
assign MEM[10120] = MEM[4517] + MEM[7516];
assign MEM[10121] = MEM[4726] + MEM[7828];
assign MEM[10122] = MEM[4770] + MEM[7529];
assign MEM[10123] = MEM[4780] + MEM[7569];
assign MEM[10124] = MEM[4783] + MEM[7532];
assign MEM[10125] = MEM[4861] + MEM[7914];
assign MEM[10126] = MEM[5139] + MEM[7968];
assign MEM[10127] = MEM[5282] + MEM[7866];
assign MEM[10128] = MEM[5315] + MEM[6079];
assign MEM[10129] = MEM[5558] + MEM[7490];
assign MEM[10130] = MEM[5754] + MEM[7812];
assign MEM[10131] = MEM[5946] + MEM[7648];
assign MEM[10132] = MEM[6195] + MEM[7630];
assign MEM[10133] = MEM[6213] + MEM[7673];
assign MEM[10134] = MEM[7260] + MEM[2023];
assign MEM[10135] = MEM[7296] + MEM[7652];
assign MEM[10136] = MEM[7399] + MEM[7629];
assign MEM[10137] = MEM[7411] + MEM[7672];
assign MEM[10138] = MEM[7418] + MEM[7674];
assign MEM[10139] = MEM[7433] + MEM[7663];
assign MEM[10140] = MEM[7436] + MEM[3802];
assign MEM[10141] = MEM[7440] + MEM[7710];
assign MEM[10142] = MEM[7448] + MEM[7683];
assign MEM[10143] = MEM[7450] + MEM[7669];
assign MEM[10144] = MEM[7453] + MEM[7617];
assign MEM[10145] = MEM[7456] + MEM[7485];
assign MEM[10146] = MEM[7463] + MEM[8013];
assign MEM[10147] = MEM[7465] + MEM[7730];
assign MEM[10148] = MEM[7484] + MEM[3006];
assign MEM[10149] = MEM[7500] + MEM[7888];
assign MEM[10150] = MEM[7559] + MEM[7677];
assign MEM[10151] = MEM[7568] + MEM[7781];
assign MEM[10152] = MEM[7577] + MEM[7656];
assign MEM[10153] = MEM[7579] + MEM[7778];
assign MEM[10154] = MEM[7581] + MEM[2663];
assign MEM[10155] = MEM[7596] + MEM[7681];
assign MEM[10156] = MEM[7608] + MEM[4958];
assign MEM[10157] = MEM[7619] + MEM[2109];
assign MEM[10158] = MEM[7624] + MEM[2620];
assign MEM[10159] = MEM[7660] + MEM[7702];
assign MEM[10160] = MEM[7670] + MEM[7709];
assign MEM[10161] = MEM[7671] + MEM[7713];
assign MEM[10162] = MEM[7675] + MEM[7632];
assign MEM[10163] = MEM[7679] + MEM[7799];
assign MEM[10164] = MEM[7686] + MEM[7718];
assign MEM[10165] = MEM[7688] + MEM[7772];
assign MEM[10166] = MEM[7691] + MEM[7788];
assign MEM[10167] = MEM[7694] + MEM[5722];
assign MEM[10168] = MEM[7699] + MEM[8431];
assign MEM[10169] = MEM[7700] + MEM[7764];
assign MEM[10170] = MEM[7712] + MEM[7857];
assign MEM[10171] = MEM[7717] + MEM[7858];
assign MEM[10172] = MEM[7729] + MEM[7986];
assign MEM[10173] = MEM[7749] + MEM[3234];
assign MEM[10174] = MEM[7758] + MEM[7820];
assign MEM[10175] = MEM[7761] + MEM[8438];
assign MEM[10176] = MEM[7762] + MEM[2527];
assign MEM[10177] = MEM[7765] + MEM[8037];
assign MEM[10178] = MEM[7773] + MEM[8136];
assign MEM[10179] = MEM[7783] + MEM[7956];
assign MEM[10180] = MEM[7792] + MEM[3183];
assign MEM[10181] = MEM[7804] + MEM[4907];
assign MEM[10182] = MEM[7810] + MEM[8208];
assign MEM[10183] = MEM[7825] + MEM[3034];
assign MEM[10184] = MEM[7840] + MEM[3502];
assign MEM[10185] = MEM[7846] + MEM[8186];
assign MEM[10186] = MEM[7850] + MEM[7915];
assign MEM[10187] = MEM[7859] + MEM[7946];
assign MEM[10188] = MEM[7863] + MEM[3771];
assign MEM[10189] = MEM[7870] + MEM[7980];
assign MEM[10190] = MEM[7874] + MEM[7926];
assign MEM[10191] = MEM[7891] + MEM[8097];
assign MEM[10192] = MEM[7897] + MEM[8141];
assign MEM[10193] = MEM[7913] + MEM[959];
assign MEM[10194] = MEM[7918] + MEM[5324];
assign MEM[10195] = MEM[7929] + MEM[7875];
assign MEM[10196] = MEM[7938] + MEM[2407];
assign MEM[10197] = MEM[7948] + MEM[7647];
assign MEM[10198] = MEM[7967] + MEM[7961];
assign MEM[10199] = MEM[7982] + MEM[8031];
assign MEM[10200] = MEM[8007] + MEM[7937];
assign MEM[10201] = MEM[8012] + MEM[4475];
assign MEM[10202] = MEM[8035] + MEM[8113];
assign MEM[10203] = MEM[8052] + MEM[8140];
assign MEM[10204] = MEM[8064] + MEM[8044];
assign MEM[10205] = MEM[8070] + MEM[8189];
assign MEM[10206] = MEM[8117] + MEM[8321];
assign MEM[10207] = MEM[8118] + MEM[8673];
assign MEM[10208] = MEM[8120] + MEM[3235];
assign MEM[10209] = MEM[8127] + MEM[8193];
assign MEM[10210] = MEM[8129] + MEM[8166];
assign MEM[10211] = MEM[8178] + MEM[7653];
assign MEM[10212] = MEM[8195] + MEM[7838];
assign MEM[10213] = MEM[8224] + MEM[8407];
assign MEM[10214] = MEM[8288] + MEM[7887];
assign MEM[10215] = MEM[8359] + MEM[8522];
assign MEM[10216] = MEM[8390] + MEM[7940];
assign MEM[10217] = MEM[8393] + MEM[8936];
assign MEM[10218] = MEM[8394] + MEM[8179];
assign MEM[10219] = MEM[8474] + MEM[7871];
assign MEM[10220] = MEM[135] + MEM[3525];
assign MEM[10221] = MEM[183] + MEM[8354];
assign MEM[10222] = MEM[382] + MEM[7685];
assign MEM[10223] = MEM[542] + MEM[2086];
assign MEM[10224] = MEM[854] + MEM[7535];
assign MEM[10225] = MEM[978] + MEM[8307];
assign MEM[10226] = MEM[1119] + MEM[2764];
assign MEM[10227] = MEM[1126] + MEM[4533];
assign MEM[10228] = MEM[1178] + MEM[8368];
assign MEM[10229] = MEM[1438] + MEM[8021];
assign MEM[10230] = MEM[1550] + MEM[7939];
assign MEM[10231] = MEM[1820] + MEM[5987];
assign MEM[10232] = MEM[2013] + MEM[8128];
assign MEM[10233] = MEM[2126] + MEM[3438];
assign MEM[10234] = MEM[2253] + MEM[3396];
assign MEM[10235] = MEM[2269] + MEM[7714];
assign MEM[10236] = MEM[2372] + MEM[7734];
assign MEM[10237] = MEM[2574] + MEM[3164];
assign MEM[10238] = MEM[2607] + MEM[5991];
assign MEM[10239] = MEM[2629] + MEM[8024];
assign MEM[10240] = MEM[2983] + MEM[7662];
assign MEM[10241] = MEM[3366] + MEM[7798];
assign MEM[10242] = MEM[3484] + MEM[7950];
assign MEM[10243] = MEM[3763] + MEM[7658];
assign MEM[10244] = MEM[3909] + MEM[7748];
assign MEM[10245] = MEM[4022] + MEM[6167];
assign MEM[10246] = MEM[4195] + MEM[5461];
assign MEM[10247] = MEM[4252] + MEM[7974];
assign MEM[10248] = MEM[4286] + MEM[7809];
assign MEM[10249] = MEM[4445] + MEM[8068];
assign MEM[10250] = MEM[4563] + MEM[7844];
assign MEM[10251] = MEM[4718] + MEM[7784];
assign MEM[10252] = MEM[4775] + MEM[7805];
assign MEM[10253] = MEM[4906] + MEM[7590];
assign MEM[10254] = MEM[5012] + MEM[7779];
assign MEM[10255] = MEM[5022] + MEM[7644];
assign MEM[10256] = MEM[5029] + MEM[8346];
assign MEM[10257] = MEM[5038] + MEM[7848];
assign MEM[10258] = MEM[5341] + MEM[5892];
assign MEM[10259] = MEM[5403] + MEM[8041];
assign MEM[10260] = MEM[5623] + MEM[7498];
assign MEM[10261] = MEM[5627] + MEM[7845];
assign MEM[10262] = MEM[5658] + MEM[8106];
assign MEM[10263] = MEM[5702] + MEM[7721];
assign MEM[10264] = MEM[6143] + MEM[7879];
assign MEM[10265] = MEM[6215] + MEM[8071];
assign MEM[10266] = MEM[7504] + MEM[8062];
assign MEM[10267] = MEM[7509] + MEM[7867];
assign MEM[10268] = MEM[7626] + MEM[7780];
assign MEM[10269] = MEM[7650] + MEM[7736];
assign MEM[10270] = MEM[7655] + MEM[8269];
assign MEM[10271] = MEM[7659] + MEM[8074];
assign MEM[10272] = MEM[7687] + MEM[7971];
assign MEM[10273] = MEM[7693] + MEM[8272];
assign MEM[10274] = MEM[7705] + MEM[7818];
assign MEM[10275] = MEM[7708] + MEM[7941];
assign MEM[10276] = MEM[7716] + MEM[8059];
assign MEM[10277] = MEM[7719] + MEM[8247];
assign MEM[10278] = MEM[7722] + MEM[7732];
assign MEM[10279] = MEM[7724] + MEM[7930];
assign MEM[10280] = MEM[7726] + MEM[7886];
assign MEM[10281] = MEM[7728] + MEM[7750];
assign MEM[10282] = MEM[7738] + MEM[8014];
assign MEM[10283] = MEM[7754] + MEM[7755];
assign MEM[10284] = MEM[7759] + MEM[7795];
assign MEM[10285] = MEM[7766] + MEM[3869];
assign MEM[10286] = MEM[7770] + MEM[2763];
assign MEM[10287] = MEM[7774] + MEM[8015];
assign MEM[10288] = MEM[7793] + MEM[7957];
assign MEM[10289] = MEM[7803] + MEM[8077];
assign MEM[10290] = MEM[7806] + MEM[7989];
assign MEM[10291] = MEM[7811] + MEM[8078];
assign MEM[10292] = MEM[7819] + MEM[301];
assign MEM[10293] = MEM[7826] + MEM[7964];
assign MEM[10294] = MEM[7835] + MEM[8018];
assign MEM[10295] = MEM[7851] + MEM[8146];
assign MEM[10296] = MEM[7861] + MEM[1188];
assign MEM[10297] = MEM[7876] + MEM[8010];
assign MEM[10298] = MEM[7877] + MEM[7959];
assign MEM[10299] = MEM[7878] + MEM[2292];
assign MEM[10300] = MEM[7880] + MEM[8268];
assign MEM[10301] = MEM[7884] + MEM[8067];
assign MEM[10302] = MEM[7889] + MEM[8000];
assign MEM[10303] = MEM[7890] + MEM[8119];
assign MEM[10304] = MEM[7900] + MEM[8320];
assign MEM[10305] = MEM[7901] + MEM[7924];
assign MEM[10306] = MEM[7902] + MEM[8003];
assign MEM[10307] = MEM[7904] + MEM[8008];
assign MEM[10308] = MEM[7908] + MEM[8038];
assign MEM[10309] = MEM[7910] + MEM[8104];
assign MEM[10310] = MEM[7911] + MEM[8397];
assign MEM[10311] = MEM[7912] + MEM[7983];
assign MEM[10312] = MEM[7922] + MEM[8225];
assign MEM[10313] = MEM[7923] + MEM[8145];
assign MEM[10314] = MEM[7925] + MEM[8173];
assign MEM[10315] = MEM[7927] + MEM[8207];
assign MEM[10316] = MEM[7931] + MEM[8168];
assign MEM[10317] = MEM[7933] + MEM[8363];
assign MEM[10318] = MEM[7942] + MEM[8518];
assign MEM[10319] = MEM[7947] + MEM[2566];
assign MEM[10320] = MEM[7949] + MEM[8585];
assign MEM[10321] = MEM[7951] + MEM[8023];
assign MEM[10322] = MEM[7952] + MEM[8180];
assign MEM[10323] = MEM[7966] + MEM[8211];
assign MEM[10324] = MEM[7969] + MEM[8199];
assign MEM[10325] = MEM[7973] + MEM[7978];
assign MEM[10326] = MEM[7977] + MEM[8176];
assign MEM[10327] = MEM[7979] + MEM[1534];
assign MEM[10328] = MEM[7981] + MEM[7903];
assign MEM[10329] = MEM[7984] + MEM[8090];
assign MEM[10330] = MEM[7992] + MEM[8513];
assign MEM[10331] = MEM[7994] + MEM[8580];
assign MEM[10332] = MEM[7999] + MEM[8004];
assign MEM[10333] = MEM[8001] + MEM[8017];
assign MEM[10334] = MEM[8006] + MEM[8355];
assign MEM[10335] = MEM[8009] + MEM[8022];
assign MEM[10336] = MEM[8016] + MEM[8046];
assign MEM[10337] = MEM[8030] + MEM[8260];
assign MEM[10338] = MEM[8032] + MEM[8262];
assign MEM[10339] = MEM[8043] + MEM[8329];
assign MEM[10340] = MEM[8054] + MEM[8348];
assign MEM[10341] = MEM[8056] + MEM[8105];
assign MEM[10342] = MEM[8057] + MEM[8296];
assign MEM[10343] = MEM[8079] + MEM[8259];
assign MEM[10344] = MEM[8081] + MEM[8182];
assign MEM[10345] = MEM[8086] + MEM[4990];
assign MEM[10346] = MEM[8087] + MEM[4927];
assign MEM[10347] = MEM[8088] + MEM[8102];
assign MEM[10348] = MEM[8089] + MEM[8664];
assign MEM[10349] = MEM[8091] + MEM[8313];
assign MEM[10350] = MEM[8096] + MEM[8115];
assign MEM[10351] = MEM[8103] + MEM[8185];
assign MEM[10352] = MEM[8110] + MEM[8667];
assign MEM[10353] = MEM[8121] + MEM[8403];
assign MEM[10354] = MEM[8125] + MEM[8400];
assign MEM[10355] = MEM[8126] + MEM[8372];
assign MEM[10356] = MEM[8130] + MEM[8250];
assign MEM[10357] = MEM[8135] + MEM[8160];
assign MEM[10358] = MEM[8137] + MEM[8310];
assign MEM[10359] = MEM[8138] + MEM[8213];
assign MEM[10360] = MEM[8139] + MEM[8174];
assign MEM[10361] = MEM[8143] + MEM[8239];
assign MEM[10362] = MEM[8144] + MEM[8387];
assign MEM[10363] = MEM[8159] + MEM[8034];
assign MEM[10364] = MEM[8161] + MEM[8305];
assign MEM[10365] = MEM[8201] + MEM[8327];
assign MEM[10366] = MEM[8209] + MEM[8256];
assign MEM[10367] = MEM[8212] + MEM[7920];
assign MEM[10368] = MEM[8214] + MEM[8392];
assign MEM[10369] = MEM[8230] + MEM[8505];
assign MEM[10370] = MEM[8254] + MEM[1983];
assign MEM[10371] = MEM[8270] + MEM[8409];
assign MEM[10372] = MEM[8275] + MEM[8061];
assign MEM[10373] = MEM[8277] + MEM[8076];
assign MEM[10374] = MEM[8278] + MEM[8065];
assign MEM[10375] = MEM[8279] + MEM[8232];
assign MEM[10376] = MEM[8292] + MEM[8124];
assign MEM[10377] = MEM[8293] + MEM[8190];
assign MEM[10378] = MEM[8300] + MEM[8384];
assign MEM[10379] = MEM[8312] + MEM[8626];
assign MEM[10380] = MEM[8317] + MEM[8674];
assign MEM[10381] = MEM[8331] + MEM[8383];
assign MEM[10382] = MEM[8332] + MEM[8050];
assign MEM[10383] = MEM[8351] + MEM[8162];
assign MEM[10384] = MEM[8378] + MEM[7932];
assign MEM[10385] = MEM[8386] + MEM[8281];
assign MEM[10386] = MEM[8388] + MEM[8682];
assign MEM[10387] = MEM[8402] + MEM[8947];
assign MEM[10388] = MEM[8405] + MEM[8642];
assign MEM[10389] = MEM[8406] + MEM[8297];
assign MEM[10390] = MEM[8410] + MEM[7767];
assign MEM[10391] = MEM[8412] + MEM[8486];
assign MEM[10392] = MEM[8502] + MEM[8316];
assign MEM[10393] = MEM[8529] + MEM[7993];
assign MEM[10394] = MEM[8549] + MEM[8072];
assign MEM[10395] = MEM[8567] + MEM[8323];
assign MEM[10396] = MEM[8608] + MEM[8657];
assign MEM[10397] = MEM[8614] + MEM[8548];
assign MEM[10398] = MEM[8658] + MEM[8733];
assign MEM[10399] = MEM[8677] + MEM[8205];
assign MEM[10400] = MEM[8678] + MEM[8546];
assign MEM[10401] = MEM[8684] + MEM[8020];
assign MEM[10402] = MEM[8696] + MEM[8645];
assign MEM[10403] = MEM[8939] + MEM[8528];
assign MEM[10404] = MEM[8950] + MEM[8715];
assign MEM[10405] = MEM[9201] + MEM[8994];
assign MEM[10406] = MEM[9203] + MEM[8426];
assign MEM[10407] = MEM[9449] + MEM[8670];
assign MEM[10408] = MEM[9466] + MEM[8873];
assign MEM[10409] = MEM[746] + MEM[8051];
assign MEM[10410] = MEM[931] + MEM[8427];
assign MEM[10411] = MEM[982] + MEM[8083];
assign MEM[10412] = MEM[1026] + MEM[8058];
assign MEM[10413] = MEM[1158] + MEM[1869];
assign MEM[10414] = MEM[1196] + MEM[8220];
assign MEM[10415] = MEM[1237] + MEM[8510];
assign MEM[10416] = MEM[1718] + MEM[7917];
assign MEM[10417] = MEM[1903] + MEM[8019];
assign MEM[10418] = MEM[2354] + MEM[8285];
assign MEM[10419] = MEM[2634] + MEM[8063];
assign MEM[10420] = MEM[2717] + MEM[8175];
assign MEM[10421] = MEM[2814] + MEM[8381];
assign MEM[10422] = MEM[3178] + MEM[8183];
assign MEM[10423] = MEM[3198] + MEM[4413];
assign MEM[10424] = MEM[3266] + MEM[8242];
assign MEM[10425] = MEM[3439] + MEM[8309];
assign MEM[10426] = MEM[4227] + MEM[9354];
assign MEM[10427] = MEM[4422] + MEM[1708];
assign MEM[10428] = MEM[4562] + MEM[4570];
assign MEM[10429] = MEM[5212] + MEM[8391];
assign MEM[10430] = MEM[5430] + MEM[8123];
assign MEM[10431] = MEM[5706] + MEM[3267];
assign MEM[10432] = MEM[5895] + MEM[8314];
assign MEM[10433] = MEM[5940] + MEM[8085];
assign MEM[10434] = MEM[6039] + MEM[8399];
assign MEM[10435] = MEM[6140] + MEM[8027];
assign MEM[10436] = MEM[6159] + MEM[8203];
assign MEM[10437] = MEM[7849] + MEM[8353];
assign MEM[10438] = MEM[7892] + MEM[8306];
assign MEM[10439] = MEM[7898] + MEM[8217];
assign MEM[10440] = MEM[7899] + MEM[8448];
assign MEM[10441] = MEM[7909] + MEM[8228];
assign MEM[10442] = MEM[7928] + MEM[8817];
assign MEM[10443] = MEM[7943] + MEM[8206];
assign MEM[10444] = MEM[7960] + MEM[8286];
assign MEM[10445] = MEM[7972] + MEM[4138];
assign MEM[10446] = MEM[7985] + MEM[8233];
assign MEM[10447] = MEM[7987] + MEM[8194];
assign MEM[10448] = MEM[7995] + MEM[8241];
assign MEM[10449] = MEM[7997] + MEM[9530];
assign MEM[10450] = MEM[8002] + MEM[8069];
assign MEM[10451] = MEM[8011] + MEM[8219];
assign MEM[10452] = MEM[8025] + MEM[8155];
assign MEM[10453] = MEM[8040] + MEM[8411];
assign MEM[10454] = MEM[8060] + MEM[996];
assign MEM[10455] = MEM[8073] + MEM[8238];
assign MEM[10456] = MEM[8075] + MEM[8165];
assign MEM[10457] = MEM[8082] + MEM[8234];
assign MEM[10458] = MEM[8099] + MEM[8417];
assign MEM[10459] = MEM[8101] + MEM[8147];
assign MEM[10460] = MEM[8111] + MEM[8325];
assign MEM[10461] = MEM[8122] + MEM[8563];
assign MEM[10462] = MEM[8142] + MEM[8164];
assign MEM[10463] = MEM[8149] + MEM[8248];
assign MEM[10464] = MEM[8163] + MEM[5766];
assign MEM[10465] = MEM[8167] + MEM[8172];
assign MEM[10466] = MEM[8170] + MEM[8229];
assign MEM[10467] = MEM[8181] + MEM[8215];
assign MEM[10468] = MEM[8187] + MEM[8227];
assign MEM[10469] = MEM[8188] + MEM[8477];
assign MEM[10470] = MEM[8200] + MEM[3516];
assign MEM[10471] = MEM[8204] + MEM[8319];
assign MEM[10472] = MEM[8210] + MEM[8338];
assign MEM[10473] = MEM[8216] + MEM[8360];
assign MEM[10474] = MEM[8221] + MEM[8290];
assign MEM[10475] = MEM[8223] + MEM[8334];
assign MEM[10476] = MEM[8236] + MEM[8496];
assign MEM[10477] = MEM[8237] + MEM[8261];
assign MEM[10478] = MEM[8244] + MEM[8834];
assign MEM[10479] = MEM[8246] + MEM[8509];
assign MEM[10480] = MEM[8249] + MEM[8251];
assign MEM[10481] = MEM[8253] + MEM[8534];
assign MEM[10482] = MEM[8255] + MEM[8471];
assign MEM[10483] = MEM[8258] + MEM[8499];
assign MEM[10484] = MEM[8263] + MEM[8443];
assign MEM[10485] = MEM[8264] + MEM[8436];
assign MEM[10486] = MEM[8265] + MEM[8532];
assign MEM[10487] = MEM[8267] + MEM[8781];
assign MEM[10488] = MEM[8280] + MEM[8301];
assign MEM[10489] = MEM[8287] + MEM[8850];
assign MEM[10490] = MEM[8289] + MEM[8704];
assign MEM[10491] = MEM[8295] + MEM[8454];
assign MEM[10492] = MEM[8298] + MEM[8515];
assign MEM[10493] = MEM[8303] + MEM[8235];
assign MEM[10494] = MEM[8304] + MEM[8690];
assign MEM[10495] = MEM[8308] + MEM[8555];
assign MEM[10496] = MEM[8311] + MEM[8243];
assign MEM[10497] = MEM[8318] + MEM[8668];
assign MEM[10498] = MEM[8326] + MEM[8597];
assign MEM[10499] = MEM[8330] + MEM[8851];
assign MEM[10500] = MEM[8335] + MEM[3830];
assign MEM[10501] = MEM[8336] + MEM[8475];
assign MEM[10502] = MEM[8340] + MEM[8646];
assign MEM[10503] = MEM[8344] + MEM[8732];
assign MEM[10504] = MEM[8347] + MEM[8369];
assign MEM[10505] = MEM[8352] + MEM[8570];
assign MEM[10506] = MEM[8356] + MEM[8564];
assign MEM[10507] = MEM[8357] + MEM[8800];
assign MEM[10508] = MEM[8358] + MEM[8881];
assign MEM[10509] = MEM[8361] + MEM[8521];
assign MEM[10510] = MEM[8362] + MEM[8790];
assign MEM[10511] = MEM[8365] + MEM[8408];
assign MEM[10512] = MEM[8367] + MEM[8492];
assign MEM[10513] = MEM[8377] + MEM[8611];
assign MEM[10514] = MEM[8380] + MEM[8530];
assign MEM[10515] = MEM[8385] + MEM[8437];
assign MEM[10516] = MEM[8389] + MEM[8418];
assign MEM[10517] = MEM[8398] + MEM[2090];
assign MEM[10518] = MEM[8401] + MEM[8192];
assign MEM[10519] = MEM[8404] + MEM[8757];
assign MEM[10520] = MEM[8429] + MEM[8907];
assign MEM[10521] = MEM[8435] + MEM[8171];
assign MEM[10522] = MEM[8444] + MEM[8899];
assign MEM[10523] = MEM[8447] + MEM[8271];
assign MEM[10524] = MEM[8455] + MEM[8550];
assign MEM[10525] = MEM[8460] + MEM[8487];
assign MEM[10526] = MEM[8463] + MEM[9217];
assign MEM[10527] = MEM[8469] + MEM[8503];
assign MEM[10528] = MEM[8478] + MEM[8531];
assign MEM[10529] = MEM[8491] + MEM[8575];
assign MEM[10530] = MEM[8494] + MEM[8276];
assign MEM[10531] = MEM[8495] + MEM[8771];
assign MEM[10532] = MEM[8504] + MEM[8562];
assign MEM[10533] = MEM[8514] + MEM[8095];
assign MEM[10534] = MEM[8527] + MEM[8432];
assign MEM[10535] = MEM[8533] + MEM[8773];
assign MEM[10536] = MEM[8542] + MEM[8766];
assign MEM[10537] = MEM[8552] + MEM[8601];
assign MEM[10538] = MEM[8558] + MEM[8579];
assign MEM[10539] = MEM[8561] + MEM[8683];
assign MEM[10540] = MEM[8573] + MEM[8364];
assign MEM[10541] = MEM[8578] + MEM[8445];
assign MEM[10542] = MEM[8589] + MEM[8282];
assign MEM[10543] = MEM[8591] + MEM[8458];
assign MEM[10544] = MEM[8599] + MEM[8675];
assign MEM[10545] = MEM[8603] + MEM[8080];
assign MEM[10546] = MEM[8605] + MEM[8456];
assign MEM[10547] = MEM[8609] + MEM[8648];
assign MEM[10548] = MEM[8619] + MEM[8654];
assign MEM[10549] = MEM[8630] + MEM[9269];
assign MEM[10550] = MEM[8638] + MEM[8291];
assign MEM[10551] = MEM[8644] + MEM[9064];
assign MEM[10552] = MEM[8655] + MEM[8931];
assign MEM[10553] = MEM[8660] + MEM[8661];
assign MEM[10554] = MEM[8666] + MEM[8695];
assign MEM[10555] = MEM[8686] + MEM[8470];
assign MEM[10556] = MEM[8687] + MEM[8745];
assign MEM[10557] = MEM[8699] + MEM[8366];
assign MEM[10558] = MEM[8723] + MEM[9104];
assign MEM[10559] = MEM[8754] + MEM[8540];
assign MEM[10560] = MEM[8768] + MEM[8938];
assign MEM[10561] = MEM[8804] + MEM[8904];
assign MEM[10562] = MEM[8839] + MEM[8997];
assign MEM[10563] = MEM[8863] + MEM[8441];
assign MEM[10564] = MEM[8910] + MEM[8672];
assign MEM[10565] = MEM[8913] + MEM[8741];
assign MEM[10566] = MEM[8921] + MEM[9213];
assign MEM[10567] = MEM[8942] + MEM[9192];
assign MEM[10568] = MEM[8944] + MEM[8940];
assign MEM[10569] = MEM[8962] + MEM[2235];
assign MEM[10570] = MEM[9020] + MEM[8595];
assign MEM[10571] = MEM[9214] + MEM[9272];
assign MEM[10572] = MEM[9373] + MEM[9051];
assign MEM[10573] = MEM[509] + MEM[8302];
assign MEM[10574] = MEM[1007] + MEM[8610];
assign MEM[10575] = MEM[1046] + MEM[8266];
assign MEM[10576] = MEM[1906] + MEM[8433];
assign MEM[10577] = MEM[3892] + MEM[1509];
assign MEM[10578] = MEM[4019] + MEM[8257];
assign MEM[10579] = MEM[4197] + MEM[8596];
assign MEM[10580] = MEM[4458] + MEM[8520];
assign MEM[10581] = MEM[4597] + MEM[8333];
assign MEM[10582] = MEM[4899] + MEM[8765];
assign MEM[10583] = MEM[5797] + MEM[8396];
assign MEM[10584] = MEM[8202] + MEM[5294];
assign MEM[10585] = MEM[8222] + MEM[8274];
assign MEM[10586] = MEM[8231] + MEM[8294];
assign MEM[10587] = MEM[8240] + MEM[8468];
assign MEM[10588] = MEM[8245] + MEM[8717];
assign MEM[10589] = MEM[8252] + MEM[8450];
assign MEM[10590] = MEM[8273] + MEM[8416];
assign MEM[10591] = MEM[8284] + MEM[8371];
assign MEM[10592] = MEM[8299] + MEM[8419];
assign MEM[10593] = MEM[8315] + MEM[8526];
assign MEM[10594] = MEM[8322] + MEM[8461];
assign MEM[10595] = MEM[8324] + MEM[8618];
assign MEM[10596] = MEM[8339] + MEM[8777];
assign MEM[10597] = MEM[8349] + MEM[8395];
assign MEM[10598] = MEM[8370] + MEM[3260];
assign MEM[10599] = MEM[8376] + MEM[8382];
assign MEM[10600] = MEM[8379] + MEM[8551];
assign MEM[10601] = MEM[8420] + MEM[8517];
assign MEM[10602] = MEM[8424] + MEM[8442];
assign MEM[10603] = MEM[8425] + MEM[8434];
assign MEM[10604] = MEM[8428] + MEM[8890];
assign MEM[10605] = MEM[8430] + MEM[8764];
assign MEM[10606] = MEM[8439] + MEM[8653];
assign MEM[10607] = MEM[8440] + MEM[8671];
assign MEM[10608] = MEM[8446] + MEM[8598];
assign MEM[10609] = MEM[8451] + MEM[8697];
assign MEM[10610] = MEM[8452] + MEM[8967];
assign MEM[10611] = MEM[8457] + MEM[8539];
assign MEM[10612] = MEM[8459] + MEM[8693];
assign MEM[10613] = MEM[8462] + MEM[8786];
assign MEM[10614] = MEM[8464] + MEM[8996];
assign MEM[10615] = MEM[8466] + MEM[8681];
assign MEM[10616] = MEM[8472] + MEM[8554];
assign MEM[10617] = MEM[8473] + MEM[8738];
assign MEM[10618] = MEM[8476] + MEM[9003];
assign MEM[10619] = MEM[8480] + MEM[8787];
assign MEM[10620] = MEM[8481] + MEM[4962];
assign MEM[10621] = MEM[8482] + MEM[9110];
assign MEM[10622] = MEM[8484] + MEM[8751];
assign MEM[10623] = MEM[8485] + MEM[9013];
assign MEM[10624] = MEM[8489] + MEM[8679];
assign MEM[10625] = MEM[8490] + MEM[8830];
assign MEM[10626] = MEM[8497] + MEM[8847];
assign MEM[10627] = MEM[8498] + MEM[8640];
assign MEM[10628] = MEM[8500] + MEM[8689];
assign MEM[10629] = MEM[8501] + MEM[8537];
assign MEM[10630] = MEM[8511] + MEM[8524];
assign MEM[10631] = MEM[8519] + MEM[8853];
assign MEM[10632] = MEM[8523] + MEM[8590];
assign MEM[10633] = MEM[8525] + MEM[8784];
assign MEM[10634] = MEM[8538] + MEM[8566];
assign MEM[10635] = MEM[8541] + MEM[8621];
assign MEM[10636] = MEM[8544] + MEM[8791];
assign MEM[10637] = MEM[8553] + MEM[8577];
assign MEM[10638] = MEM[8556] + MEM[8565];
assign MEM[10639] = MEM[8559] + MEM[8694];
assign MEM[10640] = MEM[8560] + MEM[8837];
assign MEM[10641] = MEM[8574] + MEM[8636];
assign MEM[10642] = MEM[8576] + MEM[8583];
assign MEM[10643] = MEM[8581] + MEM[8772];
assign MEM[10644] = MEM[8582] + MEM[8612];
assign MEM[10645] = MEM[8584] + MEM[8669];
assign MEM[10646] = MEM[8586] + MEM[8908];
assign MEM[10647] = MEM[8587] + MEM[9025];
assign MEM[10648] = MEM[8588] + MEM[9009];
assign MEM[10649] = MEM[8600] + MEM[8729];
assign MEM[10650] = MEM[8602] + MEM[8780];
assign MEM[10651] = MEM[8604] + MEM[8937];
assign MEM[10652] = MEM[8606] + MEM[9221];
assign MEM[10653] = MEM[8607] + MEM[8972];
assign MEM[10654] = MEM[8613] + MEM[8727];
assign MEM[10655] = MEM[8615] + MEM[9124];
assign MEM[10656] = MEM[8617] + MEM[8632];
assign MEM[10657] = MEM[8620] + MEM[8760];
assign MEM[10658] = MEM[8622] + MEM[9011];
assign MEM[10659] = MEM[8637] + MEM[8647];
assign MEM[10660] = MEM[8639] + MEM[8980];
assign MEM[10661] = MEM[8641] + MEM[8812];
assign MEM[10662] = MEM[8651] + MEM[8862];
assign MEM[10663] = MEM[8652] + MEM[9189];
assign MEM[10664] = MEM[8656] + MEM[8728];
assign MEM[10665] = MEM[8659] + MEM[8861];
assign MEM[10666] = MEM[8662] + MEM[8746];
assign MEM[10667] = MEM[8663] + MEM[8734];
assign MEM[10668] = MEM[8665] + MEM[8731];
assign MEM[10669] = MEM[8688] + MEM[8845];
assign MEM[10670] = MEM[8692] + MEM[8718];
assign MEM[10671] = MEM[8707] + MEM[8941];
assign MEM[10672] = MEM[8711] + MEM[8880];
assign MEM[10673] = MEM[8714] + MEM[9026];
assign MEM[10674] = MEM[8719] + MEM[9199];
assign MEM[10675] = MEM[8720] + MEM[8943];
assign MEM[10676] = MEM[8722] + MEM[9090];
assign MEM[10677] = MEM[8725] + MEM[8756];
assign MEM[10678] = MEM[8726] + MEM[8767];
assign MEM[10679] = MEM[8740] + MEM[9215];
assign MEM[10680] = MEM[8747] + MEM[8917];
assign MEM[10681] = MEM[8748] + MEM[8960];
assign MEM[10682] = MEM[8749] + MEM[8846];
assign MEM[10683] = MEM[8779] + MEM[8843];
assign MEM[10684] = MEM[8789] + MEM[8721];
assign MEM[10685] = MEM[8793] + MEM[2594];
assign MEM[10686] = MEM[8803] + MEM[8866];
assign MEM[10687] = MEM[8808] + MEM[8932];
assign MEM[10688] = MEM[8810] + MEM[8831];
assign MEM[10689] = MEM[8818] + MEM[9177];
assign MEM[10690] = MEM[8824] + MEM[8568];
assign MEM[10691] = MEM[8841] + MEM[9115];
assign MEM[10692] = MEM[8856] + MEM[8708];
assign MEM[10693] = MEM[8865] + MEM[9258];
assign MEM[10694] = MEM[8872] + MEM[9458];
assign MEM[10695] = MEM[8874] + MEM[8976];
assign MEM[10696] = MEM[8887] + MEM[8506];
assign MEM[10697] = MEM[8896] + MEM[9059];
assign MEM[10698] = MEM[8897] + MEM[8919];
assign MEM[10699] = MEM[8909] + MEM[8783];
assign MEM[10700] = MEM[8914] + MEM[8649];
assign MEM[10701] = MEM[8920] + MEM[8536];
assign MEM[10702] = MEM[8922] + MEM[8806];
assign MEM[10703] = MEM[8924] + MEM[9296];
assign MEM[10704] = MEM[8925] + MEM[8788];
assign MEM[10705] = MEM[8929] + MEM[9070];
assign MEM[10706] = MEM[8930] + MEM[9044];
assign MEM[10707] = MEM[8935] + MEM[9106];
assign MEM[10708] = MEM[8945] + MEM[8877];
assign MEM[10709] = MEM[8946] + MEM[8927];
assign MEM[10710] = MEM[8948] + MEM[8512];
assign MEM[10711] = MEM[8951] + MEM[9145];
assign MEM[10712] = MEM[8957] + MEM[9079];
assign MEM[10713] = MEM[8958] + MEM[9651];
assign MEM[10714] = MEM[8982] + MEM[8926];
assign MEM[10715] = MEM[9035] + MEM[9047];
assign MEM[10716] = MEM[9046] + MEM[8543];
assign MEM[10717] = MEM[9058] + MEM[8959];
assign MEM[10718] = MEM[9097] + MEM[8792];
assign MEM[10719] = MEM[9105] + MEM[8989];
assign MEM[10720] = MEM[9132] + MEM[8848];
assign MEM[10721] = MEM[9147] + MEM[8878];
assign MEM[10722] = MEM[9167] + MEM[8698];
assign MEM[10723] = MEM[9193] + MEM[9356];
assign MEM[10724] = MEM[9212] + MEM[8912];
assign MEM[10725] = MEM[9218] + MEM[8983];
assign MEM[10726] = MEM[9275] + MEM[8876];
assign MEM[10727] = MEM[9357] + MEM[9144];
assign MEM[10728] = MEM[9374] + MEM[9112];
assign MEM[10729] = MEM[9392] + MEM[9232];
assign MEM[10730] = MEM[9407] + MEM[8822];
assign MEM[10731] = MEM[9416] + MEM[9010];
assign MEM[10732] = MEM[9428] + MEM[9317];
assign MEM[10733] = MEM[9429] + MEM[9313];
assign MEM[10734] = MEM[9472] + MEM[8685];
assign MEM[10735] = MEM[9750] + MEM[8849];
assign MEM[10736] = MEM[9859] + MEM[9637];
assign MEM[10737] = MEM[654] + MEM[8735];
assign MEM[10738] = MEM[663] + MEM[9062];
assign MEM[10739] = MEM[5238] + MEM[8465];
assign MEM[10740] = MEM[8414] + MEM[8752];
assign MEM[10741] = MEM[8415] + MEM[8739];
assign MEM[10742] = MEM[8479] + MEM[8545];
assign MEM[10743] = MEM[8488] + MEM[8838];
assign MEM[10744] = MEM[8516] + MEM[8737];
assign MEM[10745] = MEM[8535] + MEM[8709];
assign MEM[10746] = MEM[8557] + MEM[8807];
assign MEM[10747] = MEM[8569] + MEM[8854];
assign MEM[10748] = MEM[8571] + MEM[8763];
assign MEM[10749] = MEM[8572] + MEM[8769];
assign MEM[10750] = MEM[8616] + MEM[8676];
assign MEM[10751] = MEM[8631] + MEM[8829];
assign MEM[10752] = MEM[8643] + MEM[8744];
assign MEM[10753] = MEM[8691] + MEM[8700];
assign MEM[10754] = MEM[8705] + MEM[8724];
assign MEM[10755] = MEM[8706] + MEM[9002];
assign MEM[10756] = MEM[8710] + MEM[8761];
assign MEM[10757] = MEM[8712] + MEM[9114];
assign MEM[10758] = MEM[8713] + MEM[8805];
assign MEM[10759] = MEM[8716] + MEM[9139];
assign MEM[10760] = MEM[8730] + MEM[9032];
assign MEM[10761] = MEM[8736] + MEM[8882];
assign MEM[10762] = MEM[8742] + MEM[8911];
assign MEM[10763] = MEM[8743] + MEM[8860];
assign MEM[10764] = MEM[8750] + MEM[9172];
assign MEM[10765] = MEM[8753] + MEM[8785];
assign MEM[10766] = MEM[8755] + MEM[8801];
assign MEM[10767] = MEM[8758] + MEM[9076];
assign MEM[10768] = MEM[8762] + MEM[8905];
assign MEM[10769] = MEM[8770] + MEM[9001];
assign MEM[10770] = MEM[8775] + MEM[8956];
assign MEM[10771] = MEM[8778] + MEM[8782];
assign MEM[10772] = MEM[8795] + MEM[8859];
assign MEM[10773] = MEM[8796] + MEM[8928];
assign MEM[10774] = MEM[8797] + MEM[8970];
assign MEM[10775] = MEM[8798] + MEM[8857];
assign MEM[10776] = MEM[8799] + MEM[9023];
assign MEM[10777] = MEM[8811] + MEM[8901];
assign MEM[10778] = MEM[8816] + MEM[8844];
assign MEM[10779] = MEM[8819] + MEM[5005];
assign MEM[10780] = MEM[8820] + MEM[8891];
assign MEM[10781] = MEM[8827] + MEM[8954];
assign MEM[10782] = MEM[8828] + MEM[9235];
assign MEM[10783] = MEM[8832] + MEM[9100];
assign MEM[10784] = MEM[8833] + MEM[8879];
assign MEM[10785] = MEM[8835] + MEM[9219];
assign MEM[10786] = MEM[8842] + MEM[9175];
assign MEM[10787] = MEM[8852] + MEM[8864];
assign MEM[10788] = MEM[8858] + MEM[8999];
assign MEM[10789] = MEM[8870] + MEM[8955];
assign MEM[10790] = MEM[8871] + MEM[8963];
assign MEM[10791] = MEM[8883] + MEM[9078];
assign MEM[10792] = MEM[8884] + MEM[9169];
assign MEM[10793] = MEM[8885] + MEM[9204];
assign MEM[10794] = MEM[8886] + MEM[8953];
assign MEM[10795] = MEM[8889] + MEM[9151];
assign MEM[10796] = MEM[8892] + MEM[9021];
assign MEM[10797] = MEM[8898] + MEM[9048];
assign MEM[10798] = MEM[8900] + MEM[9314];
assign MEM[10799] = MEM[8903] + MEM[9205];
assign MEM[10800] = MEM[8906] + MEM[8915];
assign MEM[10801] = MEM[8916] + MEM[9066];
assign MEM[10802] = MEM[8918] + MEM[8952];
assign MEM[10803] = MEM[8923] + MEM[9039];
assign MEM[10804] = MEM[8933] + MEM[9063];
assign MEM[10805] = MEM[8949] + MEM[9586];
assign MEM[10806] = MEM[8968] + MEM[9057];
assign MEM[10807] = MEM[8971] + MEM[9223];
assign MEM[10808] = MEM[8973] + MEM[8998];
assign MEM[10809] = MEM[8974] + MEM[9095];
assign MEM[10810] = MEM[8975] + MEM[9295];
assign MEM[10811] = MEM[8979] + MEM[9083];
assign MEM[10812] = MEM[8981] + MEM[9149];
assign MEM[10813] = MEM[8984] + MEM[9174];
assign MEM[10814] = MEM[8985] + MEM[9073];
assign MEM[10815] = MEM[8990] + MEM[9457];
assign MEM[10816] = MEM[9004] + MEM[9061];
assign MEM[10817] = MEM[9012] + MEM[9208];
assign MEM[10818] = MEM[9014] + MEM[9168];
assign MEM[10819] = MEM[9017] + MEM[9129];
assign MEM[10820] = MEM[9018] + MEM[9122];
assign MEM[10821] = MEM[9022] + MEM[9173];
assign MEM[10822] = MEM[9027] + MEM[9016];
assign MEM[10823] = MEM[9030] + MEM[9202];
assign MEM[10824] = MEM[9033] + MEM[9138];
assign MEM[10825] = MEM[9036] + MEM[9196];
assign MEM[10826] = MEM[9045] + MEM[9242];
assign MEM[10827] = MEM[9053] + MEM[9312];
assign MEM[10828] = MEM[9054] + MEM[9360];
assign MEM[10829] = MEM[9060] + MEM[9424];
assign MEM[10830] = MEM[9080] + MEM[8802];
assign MEM[10831] = MEM[9081] + MEM[9143];
assign MEM[10832] = MEM[9082] + MEM[9395];
assign MEM[10833] = MEM[9084] + MEM[9211];
assign MEM[10834] = MEM[9089] + MEM[9195];
assign MEM[10835] = MEM[9091] + MEM[9096];
assign MEM[10836] = MEM[9092] + MEM[9140];
assign MEM[10837] = MEM[9101] + MEM[9316];
assign MEM[10838] = MEM[9108] + MEM[9085];
assign MEM[10839] = MEM[9116] + MEM[9298];
assign MEM[10840] = MEM[9118] + MEM[9234];
assign MEM[10841] = MEM[9126] + MEM[9134];
assign MEM[10842] = MEM[9130] + MEM[9233];
assign MEM[10843] = MEM[9131] + MEM[9263];
assign MEM[10844] = MEM[9136] + MEM[9606];
assign MEM[10845] = MEM[9141] + MEM[9408];
assign MEM[10846] = MEM[9146] + MEM[9262];
assign MEM[10847] = MEM[9156] + MEM[9031];
assign MEM[10848] = MEM[9157] + MEM[9093];
assign MEM[10849] = MEM[9160] + MEM[9391];
assign MEM[10850] = MEM[9166] + MEM[9150];
assign MEM[10851] = MEM[9170] + MEM[9260];
assign MEM[10852] = MEM[9176] + MEM[9318];
assign MEM[10853] = MEM[9190] + MEM[9643];
assign MEM[10854] = MEM[9197] + MEM[9207];
assign MEM[10855] = MEM[9200] + MEM[9460];
assign MEM[10856] = MEM[9206] + MEM[9338];
assign MEM[10857] = MEM[9209] + MEM[9615];
assign MEM[10858] = MEM[9220] + MEM[9111];
assign MEM[10859] = MEM[9248] + MEM[9359];
assign MEM[10860] = MEM[9250] + MEM[9152];
assign MEM[10861] = MEM[9279] + MEM[9624];
assign MEM[10862] = MEM[9284] + MEM[9321];
assign MEM[10863] = MEM[9303] + MEM[9394];
assign MEM[10864] = MEM[9331] + MEM[9447];
assign MEM[10865] = MEM[9333] + MEM[9533];
assign MEM[10866] = MEM[9337] + MEM[9024];
assign MEM[10867] = MEM[9382] + MEM[9483];
assign MEM[10868] = MEM[9399] + MEM[9075];
assign MEM[10869] = MEM[9403] + MEM[9461];
assign MEM[10870] = MEM[9409] + MEM[9431];
assign MEM[10871] = MEM[9415] + MEM[9237];
assign MEM[10872] = MEM[9437] + MEM[9326];
assign MEM[10873] = MEM[9445] + MEM[9554];
assign MEM[10874] = MEM[9455] + MEM[9297];
assign MEM[10875] = MEM[9467] + MEM[9128];
assign MEM[10876] = MEM[9468] + MEM[8823];
assign MEM[10877] = MEM[9469] + MEM[9576];
assign MEM[10878] = MEM[9470] + MEM[9664];
assign MEM[10879] = MEM[9495] + MEM[9349];
assign MEM[10880] = MEM[9535] + MEM[9266];
assign MEM[10881] = MEM[9550] + MEM[9222];
assign MEM[10882] = MEM[9557] + MEM[8987];
assign MEM[10883] = MEM[9640] + MEM[9587];
assign MEM[10884] = MEM[9641] + MEM[9121];
assign MEM[10885] = MEM[9853] + MEM[9464];
assign MEM[10886] = MEM[9862] + MEM[9538];
assign MEM[10887] = MEM[749] + MEM[9501];
assign MEM[10888] = MEM[1322] + MEM[9216];
assign MEM[10889] = MEM[3606] + MEM[9385];
assign MEM[10890] = MEM[4010] + MEM[9224];
assign MEM[10891] = MEM[4893] + MEM[8888];
assign MEM[10892] = MEM[5629] + MEM[9253];
assign MEM[10893] = MEM[8759] + MEM[9086];
assign MEM[10894] = MEM[8774] + MEM[8995];
assign MEM[10895] = MEM[8836] + MEM[9056];
assign MEM[10896] = MEM[8875] + MEM[9049];
assign MEM[10897] = MEM[8902] + MEM[8986];
assign MEM[10898] = MEM[8934] + MEM[8961];
assign MEM[10899] = MEM[8969] + MEM[9005];
assign MEM[10900] = MEM[8977] + MEM[8978];
assign MEM[10901] = MEM[8988] + MEM[9324];
assign MEM[10902] = MEM[8991] + MEM[9072];
assign MEM[10903] = MEM[8992] + MEM[9355];
assign MEM[10904] = MEM[8993] + MEM[9380];
assign MEM[10905] = MEM[9000] + MEM[9142];
assign MEM[10906] = MEM[9006] + MEM[9127];
assign MEM[10907] = MEM[9007] + MEM[9120];
assign MEM[10908] = MEM[9008] + MEM[9041];
assign MEM[10909] = MEM[9015] + MEM[9050];
assign MEM[10910] = MEM[9019] + MEM[9099];
assign MEM[10911] = MEM[9028] + MEM[9182];
assign MEM[10912] = MEM[9029] + MEM[9155];
assign MEM[10913] = MEM[9037] + MEM[9071];
assign MEM[10914] = MEM[9038] + MEM[9179];
assign MEM[10915] = MEM[9042] + MEM[9388];
assign MEM[10916] = MEM[9043] + MEM[9293];
assign MEM[10917] = MEM[9052] + MEM[9277];
assign MEM[10918] = MEM[9055] + MEM[9246];
assign MEM[10919] = MEM[9065] + MEM[9069];
assign MEM[10920] = MEM[9067] + MEM[9187];
assign MEM[10921] = MEM[9068] + MEM[9077];
assign MEM[10922] = MEM[9074] + MEM[9270];
assign MEM[10923] = MEM[9087] + MEM[9397];
assign MEM[10924] = MEM[9088] + MEM[9562];
assign MEM[10925] = MEM[9094] + MEM[9117];
assign MEM[10926] = MEM[9098] + MEM[9125];
assign MEM[10927] = MEM[9102] + MEM[9153];
assign MEM[10928] = MEM[9103] + MEM[9310];
assign MEM[10929] = MEM[9107] + MEM[9430];
assign MEM[10930] = MEM[9109] + MEM[9236];
assign MEM[10931] = MEM[9113] + MEM[9299];
assign MEM[10932] = MEM[9119] + MEM[9186];
assign MEM[10933] = MEM[9123] + MEM[9137];
assign MEM[10934] = MEM[9133] + MEM[9188];
assign MEM[10935] = MEM[9148] + MEM[9161];
assign MEM[10936] = MEM[9154] + MEM[9230];
assign MEM[10937] = MEM[9158] + MEM[9165];
assign MEM[10938] = MEM[9159] + MEM[9245];
assign MEM[10939] = MEM[9171] + MEM[9323];
assign MEM[10940] = MEM[9180] + MEM[9271];
assign MEM[10941] = MEM[9181] + MEM[9283];
assign MEM[10942] = MEM[9183] + MEM[9353];
assign MEM[10943] = MEM[9185] + MEM[9292];
assign MEM[10944] = MEM[9191] + MEM[9724];
assign MEM[10945] = MEM[9194] + MEM[9334];
assign MEM[10946] = MEM[9210] + MEM[9273];
assign MEM[10947] = MEM[9238] + MEM[9490];
assign MEM[10948] = MEM[9239] + MEM[9432];
assign MEM[10949] = MEM[9249] + MEM[9259];
assign MEM[10950] = MEM[9251] + MEM[9329];
assign MEM[10951] = MEM[9252] + MEM[9302];
assign MEM[10952] = MEM[9254] + MEM[9366];
assign MEM[10953] = MEM[9255] + MEM[9644];
assign MEM[10954] = MEM[9257] + MEM[9336];
assign MEM[10955] = MEM[9264] + MEM[9404];
assign MEM[10956] = MEM[9268] + MEM[9434];
assign MEM[10957] = MEM[9274] + MEM[9368];
assign MEM[10958] = MEM[9280] + MEM[9328];
assign MEM[10959] = MEM[9281] + MEM[9742];
assign MEM[10960] = MEM[9288] + MEM[9436];
assign MEM[10961] = MEM[9290] + MEM[9536];
assign MEM[10962] = MEM[9291] + MEM[9386];
assign MEM[10963] = MEM[9300] + MEM[9261];
assign MEM[10964] = MEM[9304] + MEM[9335];
assign MEM[10965] = MEM[9305] + MEM[319];
assign MEM[10966] = MEM[9306] + MEM[9363];
assign MEM[10967] = MEM[9307] + MEM[9352];
assign MEM[10968] = MEM[9309] + MEM[9595];
assign MEM[10969] = MEM[9319] + MEM[9320];
assign MEM[10970] = MEM[9325] + MEM[9571];
assign MEM[10971] = MEM[9327] + MEM[9514];
assign MEM[10972] = MEM[9330] + MEM[9783];
assign MEM[10973] = MEM[9341] + MEM[9528];
assign MEM[10974] = MEM[9342] + MEM[9441];
assign MEM[10975] = MEM[9343] + MEM[9267];
assign MEM[10976] = MEM[9345] + MEM[9377];
assign MEM[10977] = MEM[9348] + MEM[9362];
assign MEM[10978] = MEM[9358] + MEM[9402];
assign MEM[10979] = MEM[9375] + MEM[9425];
assign MEM[10980] = MEM[9376] + MEM[9448];
assign MEM[10981] = MEM[9381] + MEM[9390];
assign MEM[10982] = MEM[9383] + MEM[9540];
assign MEM[10983] = MEM[9384] + MEM[9655];
assign MEM[10984] = MEM[9387] + MEM[9547];
assign MEM[10985] = MEM[9401] + MEM[9301];
assign MEM[10986] = MEM[9410] + MEM[9700];
assign MEM[10987] = MEM[9413] + MEM[9607];
assign MEM[10988] = MEM[9420] + MEM[9599];
assign MEM[10989] = MEM[9421] + MEM[9657];
assign MEM[10990] = MEM[9438] + MEM[9289];
assign MEM[10991] = MEM[9443] + MEM[9364];
assign MEM[10992] = MEM[9446] + MEM[9546];
assign MEM[10993] = MEM[9451] + MEM[9600];
assign MEM[10994] = MEM[9452] + MEM[9627];
assign MEM[10995] = MEM[9454] + MEM[10125];
assign MEM[10996] = MEM[9456] + MEM[9512];
assign MEM[10997] = MEM[9474] + MEM[9620];
assign MEM[10998] = MEM[9480] + MEM[9504];
assign MEM[10999] = MEM[9487] + MEM[9244];
assign MEM[11000] = MEM[9496] + MEM[9389];
assign MEM[11001] = MEM[9502] + MEM[9583];
assign MEM[11002] = MEM[9506] + MEM[9418];
assign MEM[11003] = MEM[9508] + MEM[9597];
assign MEM[11004] = MEM[9511] + MEM[9716];
assign MEM[11005] = MEM[9513] + MEM[9560];
assign MEM[11006] = MEM[9529] + MEM[9598];
assign MEM[11007] = MEM[9539] + MEM[9498];
assign MEM[11008] = MEM[9541] + MEM[9860];
assign MEM[11009] = MEM[9542] + MEM[9713];
assign MEM[11010] = MEM[9558] + MEM[9365];
assign MEM[11011] = MEM[9569] + MEM[9656];
assign MEM[11012] = MEM[9580] + MEM[9405];
assign MEM[11013] = MEM[9588] + MEM[9198];
assign MEM[11014] = MEM[9618] + MEM[9340];
assign MEM[11015] = MEM[9623] + MEM[9427];
assign MEM[11016] = MEM[9633] + MEM[9479];
assign MEM[11017] = MEM[9635] + MEM[9393];
assign MEM[11018] = MEM[9638] + MEM[9379];
assign MEM[11019] = MEM[9647] + MEM[9505];
assign MEM[11020] = MEM[9650] + MEM[9866];
assign MEM[11021] = MEM[9654] + MEM[9619];
assign MEM[11022] = MEM[9658] + MEM[9663];
assign MEM[11023] = MEM[9671] + MEM[9412];
assign MEM[11024] = MEM[9673] + MEM[9705];
assign MEM[11025] = MEM[9675] + MEM[9577];
assign MEM[11026] = MEM[9698] + MEM[9414];
assign MEM[11027] = MEM[9712] + MEM[9423];
assign MEM[11028] = MEM[9714] + MEM[9564];
assign MEM[11029] = MEM[9735] + MEM[9520];
assign MEM[11030] = MEM[9741] + MEM[9256];
assign MEM[11031] = MEM[9758] + MEM[9411];
assign MEM[11032] = MEM[9851] + MEM[9722];
assign MEM[11033] = MEM[9981] + MEM[9034];
assign MEM[11034] = MEM[10001] + MEM[9801];
assign MEM[11035] = MEM[10173] + MEM[9994];
assign MEM[11036] = MEM[1549] + MEM[10292];
assign MEM[11037] = MEM[9178] + MEM[9509];
assign MEM[11038] = MEM[9184] + MEM[9229];
assign MEM[11039] = MEM[9228] + MEM[9243];
assign MEM[11040] = MEM[9231] + MEM[9459];
assign MEM[11041] = MEM[9240] + MEM[9282];
assign MEM[11042] = MEM[9241] + MEM[9396];
assign MEM[11043] = MEM[9247] + MEM[9351];
assign MEM[11044] = MEM[9265] + MEM[9311];
assign MEM[11045] = MEM[9276] + MEM[9625];
assign MEM[11046] = MEM[9278] + MEM[9400];
assign MEM[11047] = MEM[9285] + MEM[9473];
assign MEM[11048] = MEM[9286] + MEM[9332];
assign MEM[11049] = MEM[9287] + MEM[9372];
assign MEM[11050] = MEM[9294] + MEM[9573];
assign MEM[11051] = MEM[9308] + MEM[9476];
assign MEM[11052] = MEM[9315] + MEM[9361];
assign MEM[11053] = MEM[9322] + MEM[9440];
assign MEM[11054] = MEM[9339] + MEM[9692];
assign MEM[11055] = MEM[9344] + MEM[9485];
assign MEM[11056] = MEM[9346] + MEM[9371];
assign MEM[11057] = MEM[9347] + MEM[9350];
assign MEM[11058] = MEM[9367] + MEM[9561];
assign MEM[11059] = MEM[9369] + MEM[9515];
assign MEM[11060] = MEM[9370] + MEM[9477];
assign MEM[11061] = MEM[9378] + MEM[9559];
assign MEM[11062] = MEM[9398] + MEM[9463];
assign MEM[11063] = MEM[9406] + MEM[9422];
assign MEM[11064] = MEM[9417] + MEM[9646];
assign MEM[11065] = MEM[9419] + MEM[9521];
assign MEM[11066] = MEM[9426] + MEM[9649];
assign MEM[11067] = MEM[9433] + MEM[9453];
assign MEM[11068] = MEM[9435] + MEM[9549];
assign MEM[11069] = MEM[9439] + MEM[9450];
assign MEM[11070] = MEM[9442] + MEM[9462];
assign MEM[11071] = MEM[9444] + MEM[9652];
assign MEM[11072] = MEM[9465] + MEM[9493];
assign MEM[11073] = MEM[9471] + MEM[9747];
assign MEM[11074] = MEM[9475] + MEM[9478];
assign MEM[11075] = MEM[9481] + MEM[9829];
assign MEM[11076] = MEM[9482] + MEM[9729];
assign MEM[11077] = MEM[9484] + MEM[9737];
assign MEM[11078] = MEM[9488] + MEM[9486];
assign MEM[11079] = MEM[9489] + MEM[9537];
assign MEM[11080] = MEM[9491] + MEM[9608];
assign MEM[11081] = MEM[9494] + MEM[9567];
assign MEM[11082] = MEM[9499] + MEM[9846];
assign MEM[11083] = MEM[9503] + MEM[5919];
assign MEM[11084] = MEM[9510] + MEM[9734];
assign MEM[11085] = MEM[9516] + MEM[9621];
assign MEM[11086] = MEM[9517] + MEM[9534];
assign MEM[11087] = MEM[9518] + MEM[9695];
assign MEM[11088] = MEM[9519] + MEM[9563];
assign MEM[11089] = MEM[9522] + MEM[9578];
assign MEM[11090] = MEM[9523] + MEM[9497];
assign MEM[11091] = MEM[9524] + MEM[9631];
assign MEM[11092] = MEM[9525] + MEM[9565];
assign MEM[11093] = MEM[9526] + MEM[9531];
assign MEM[11094] = MEM[9527] + MEM[9662];
assign MEM[11095] = MEM[9532] + MEM[9822];
assign MEM[11096] = MEM[9544] + MEM[9616];
assign MEM[11097] = MEM[9545] + MEM[9548];
assign MEM[11098] = MEM[9551] + MEM[9690];
assign MEM[11099] = MEM[9552] + MEM[9957];
assign MEM[11100] = MEM[9553] + MEM[9679];
assign MEM[11101] = MEM[9555] + MEM[10010];
assign MEM[11102] = MEM[9566] + MEM[9816];
assign MEM[11103] = MEM[9568] + MEM[9761];
assign MEM[11104] = MEM[9570] + MEM[9601];
assign MEM[11105] = MEM[9572] + MEM[9574];
assign MEM[11106] = MEM[9575] + MEM[9605];
assign MEM[11107] = MEM[9579] + MEM[9592];
assign MEM[11108] = MEM[9581] + MEM[9639];
assign MEM[11109] = MEM[9584] + MEM[9794];
assign MEM[11110] = MEM[9585] + MEM[9744];
assign MEM[11111] = MEM[9589] + MEM[4750];
assign MEM[11112] = MEM[9590] + MEM[9799];
assign MEM[11113] = MEM[9591] + MEM[9766];
assign MEM[11114] = MEM[9594] + MEM[9667];
assign MEM[11115] = MEM[9596] + MEM[9720];
assign MEM[11116] = MEM[9602] + MEM[10014];
assign MEM[11117] = MEM[9603] + MEM[9790];
assign MEM[11118] = MEM[9611] + MEM[9756];
assign MEM[11119] = MEM[9613] + MEM[9719];
assign MEM[11120] = MEM[9622] + MEM[9779];
assign MEM[11121] = MEM[9626] + MEM[9838];
assign MEM[11122] = MEM[9630] + MEM[9636];
assign MEM[11123] = MEM[9632] + MEM[9802];
assign MEM[11124] = MEM[9634] + MEM[9770];
assign MEM[11125] = MEM[9642] + MEM[9686];
assign MEM[11126] = MEM[9645] + MEM[9709];
assign MEM[11127] = MEM[9660] + MEM[9681];
assign MEM[11128] = MEM[9661] + MEM[10004];
assign MEM[11129] = MEM[9665] + MEM[9971];
assign MEM[11130] = MEM[9669] + MEM[9824];
assign MEM[11131] = MEM[9688] + MEM[10017];
assign MEM[11132] = MEM[9693] + MEM[9507];
assign MEM[11133] = MEM[9702] + MEM[9668];
assign MEM[11134] = MEM[9711] + MEM[10187];
assign MEM[11135] = MEM[9717] + MEM[9803];
assign MEM[11136] = MEM[9725] + MEM[9831];
assign MEM[11137] = MEM[9727] + MEM[9894];
assign MEM[11138] = MEM[9733] + MEM[9833];
assign MEM[11139] = MEM[9738] + MEM[9707];
assign MEM[11140] = MEM[9740] + MEM[9629];
assign MEM[11141] = MEM[9746] + MEM[9847];
assign MEM[11142] = MEM[9748] + MEM[10140];
assign MEM[11143] = MEM[9762] + MEM[9823];
assign MEM[11144] = MEM[9774] + MEM[10130];
assign MEM[11145] = MEM[9780] + MEM[9969];
assign MEM[11146] = MEM[9782] + MEM[9976];
assign MEM[11147] = MEM[9791] + MEM[9844];
assign MEM[11148] = MEM[9792] + MEM[9964];
assign MEM[11149] = MEM[9796] + MEM[10052];
assign MEM[11150] = MEM[9804] + MEM[9763];
assign MEM[11151] = MEM[9808] + MEM[9967];
assign MEM[11152] = MEM[9809] + MEM[5276];
assign MEM[11153] = MEM[9817] + MEM[9870];
assign MEM[11154] = MEM[9820] + MEM[9778];
assign MEM[11155] = MEM[9830] + MEM[10101];
assign MEM[11156] = MEM[9834] + MEM[9871];
assign MEM[11157] = MEM[9839] + MEM[9730];
assign MEM[11158] = MEM[9852] + MEM[10045];
assign MEM[11159] = MEM[9855] + MEM[9896];
assign MEM[11160] = MEM[9856] + MEM[9556];
assign MEM[11161] = MEM[9864] + MEM[9899];
assign MEM[11162] = MEM[9865] + MEM[9703];
assign MEM[11163] = MEM[9872] + MEM[9906];
assign MEM[11164] = MEM[9901] + MEM[9811];
assign MEM[11165] = MEM[9912] + MEM[9953];
assign MEM[11166] = MEM[9930] + MEM[9821];
assign MEM[11167] = MEM[9985] + MEM[9492];
assign MEM[11168] = MEM[9997] + MEM[10057];
assign MEM[11169] = MEM[10032] + MEM[9875];
assign MEM[11170] = MEM[10033] + MEM[9850];
assign MEM[11171] = MEM[10035] + MEM[9781];
assign MEM[11172] = MEM[10055] + MEM[9843];
assign MEM[11173] = MEM[10058] + MEM[9837];
assign MEM[11174] = MEM[10069] + MEM[994];
assign MEM[11175] = MEM[10109] + MEM[9848];
assign MEM[11176] = MEM[10122] + MEM[9617];
assign MEM[11177] = MEM[10163] + MEM[9732];
assign MEM[11178] = MEM[847] + MEM[9827];
assign MEM[11179] = MEM[2746] + MEM[7604];
assign MEM[11180] = MEM[6575] + MEM[3274];
assign MEM[11181] = MEM[6840] + MEM[8808];
assign MEM[11182] = MEM[7002] + MEM[9897];
assign MEM[11183] = MEM[9500] + MEM[9773];
assign MEM[11184] = MEM[9543] + MEM[9697];
assign MEM[11185] = MEM[9582] + MEM[9983];
assign MEM[11186] = MEM[9593] + MEM[9836];
assign MEM[11187] = MEM[9604] + MEM[9797];
assign MEM[11188] = MEM[9609] + MEM[9689];
assign MEM[11189] = MEM[9610] + MEM[5637];
assign MEM[11190] = MEM[9612] + MEM[9683];
assign MEM[11191] = MEM[9614] + MEM[9728];
assign MEM[11192] = MEM[9628] + MEM[9788];
assign MEM[11193] = MEM[9648] + MEM[9687];
assign MEM[11194] = MEM[9653] + MEM[9682];
assign MEM[11195] = MEM[9659] + MEM[9785];
assign MEM[11196] = MEM[9666] + MEM[9826];
assign MEM[11197] = MEM[9670] + MEM[9921];
assign MEM[11198] = MEM[9672] + MEM[9752];
assign MEM[11199] = MEM[9674] + MEM[9878];
assign MEM[11200] = MEM[9677] + MEM[7509];
assign MEM[11201] = MEM[9678] + MEM[7143];
assign MEM[11202] = MEM[9680] + MEM[9694];
assign MEM[11203] = MEM[9684] + MEM[10213];
assign MEM[11204] = MEM[9685] + MEM[9793];
assign MEM[11205] = MEM[9691] + MEM[9751];
assign MEM[11206] = MEM[9696] + MEM[9753];
assign MEM[11207] = MEM[9699] + MEM[9900];
assign MEM[11208] = MEM[9704] + MEM[5461];
assign MEM[11209] = MEM[9708] + MEM[9939];
assign MEM[11210] = MEM[9710] + MEM[2507];
assign MEM[11211] = MEM[9715] + MEM[4838];
assign MEM[11212] = MEM[9718] + MEM[9755];
assign MEM[11213] = MEM[9721] + MEM[9812];
assign MEM[11214] = MEM[9723] + MEM[9828];
assign MEM[11215] = MEM[9726] + MEM[9990];
assign MEM[11216] = MEM[9731] + MEM[8274];
assign MEM[11217] = MEM[9739] + MEM[9963];
assign MEM[11218] = MEM[9743] + MEM[10070];
assign MEM[11219] = MEM[9745] + MEM[9858];
assign MEM[11220] = MEM[9749] + MEM[9992];
assign MEM[11221] = MEM[9754] + MEM[9909];
assign MEM[11222] = MEM[9757] + MEM[9941];
assign MEM[11223] = MEM[9759] + MEM[10059];
assign MEM[11224] = MEM[9760] + MEM[9892];
assign MEM[11225] = MEM[9764] + MEM[9910];
assign MEM[11226] = MEM[9765] + MEM[9810];
assign MEM[11227] = MEM[9767] + MEM[9795];
assign MEM[11228] = MEM[9768] + MEM[5780];
assign MEM[11229] = MEM[9769] + MEM[9815];
assign MEM[11230] = MEM[9771] + MEM[9922];
assign MEM[11231] = MEM[9772] + MEM[9854];
assign MEM[11232] = MEM[9775] + MEM[9789];
assign MEM[11233] = MEM[9776] + MEM[9841];
assign MEM[11234] = MEM[9777] + MEM[1799];
assign MEM[11235] = MEM[9787] + MEM[10022];
assign MEM[11236] = MEM[9798] + MEM[9807];
assign MEM[11237] = MEM[9800] + MEM[9978];
assign MEM[11238] = MEM[9805] + MEM[10247];
assign MEM[11239] = MEM[9806] + MEM[9965];
assign MEM[11240] = MEM[9813] + MEM[9880];
assign MEM[11241] = MEM[9814] + MEM[9918];
assign MEM[11242] = MEM[9818] + MEM[9885];
assign MEM[11243] = MEM[9819] + MEM[766];
assign MEM[11244] = MEM[9835] + MEM[9849];
assign MEM[11245] = MEM[9840] + MEM[3410];
assign MEM[11246] = MEM[9842] + MEM[9914];
assign MEM[11247] = MEM[9845] + MEM[5259];
assign MEM[11248] = MEM[9863] + MEM[9998];
assign MEM[11249] = MEM[9868] + MEM[10002];
assign MEM[11250] = MEM[9869] + MEM[9979];
assign MEM[11251] = MEM[9874] + MEM[9903];
assign MEM[11252] = MEM[9876] + MEM[9923];
assign MEM[11253] = MEM[9877] + MEM[10330];
assign MEM[11254] = MEM[9881] + MEM[10083];
assign MEM[11255] = MEM[9884] + MEM[9938];
assign MEM[11256] = MEM[9886] + MEM[9891];
assign MEM[11257] = MEM[9887] + MEM[9949];
assign MEM[11258] = MEM[9888] + MEM[9934];
assign MEM[11259] = MEM[9890] + MEM[9977];
assign MEM[11260] = MEM[9893] + MEM[10050];
assign MEM[11261] = MEM[9895] + MEM[10197];
assign MEM[11262] = MEM[9898] + MEM[10068];
assign MEM[11263] = MEM[9902] + MEM[540];
assign MEM[11264] = MEM[9904] + MEM[9950];
assign MEM[11265] = MEM[9905] + MEM[10020];
assign MEM[11266] = MEM[9911] + MEM[9920];
assign MEM[11267] = MEM[9913] + MEM[10179];
assign MEM[11268] = MEM[9916] + MEM[9974];
assign MEM[11269] = MEM[9917] + MEM[10000];
assign MEM[11270] = MEM[9924] + MEM[9873];
assign MEM[11271] = MEM[9925] + MEM[8002];
assign MEM[11272] = MEM[9926] + MEM[4525];
assign MEM[11273] = MEM[9928] + MEM[6141];
assign MEM[11274] = MEM[9929] + MEM[9982];
assign MEM[11275] = MEM[9932] + MEM[10018];
assign MEM[11276] = MEM[9933] + MEM[9987];
assign MEM[11277] = MEM[9935] + MEM[9947];
assign MEM[11278] = MEM[9936] + MEM[9993];
assign MEM[11279] = MEM[9937] + MEM[10123];
assign MEM[11280] = MEM[9942] + MEM[10009];
assign MEM[11281] = MEM[9944] + MEM[10030];
assign MEM[11282] = MEM[9945] + MEM[10046];
assign MEM[11283] = MEM[9946] + MEM[9706];
assign MEM[11284] = MEM[9954] + MEM[1435];
assign MEM[11285] = MEM[9959] + MEM[4309];
assign MEM[11286] = MEM[9961] + MEM[10089];
assign MEM[11287] = MEM[9962] + MEM[10023];
assign MEM[11288] = MEM[9966] + MEM[10379];
assign MEM[11289] = MEM[9968] + MEM[9786];
assign MEM[11290] = MEM[9975] + MEM[6740];
assign MEM[11291] = MEM[9986] + MEM[7848];
assign MEM[11292] = MEM[9991] + MEM[10128];
assign MEM[11293] = MEM[9996] + MEM[10201];
assign MEM[11294] = MEM[9999] + MEM[10149];
assign MEM[11295] = MEM[10003] + MEM[10162];
assign MEM[11296] = MEM[10005] + MEM[9867];
assign MEM[11297] = MEM[10007] + MEM[10177];
assign MEM[11298] = MEM[10008] + MEM[9931];
assign MEM[11299] = MEM[10019] + MEM[10147];
assign MEM[11300] = MEM[10026] + MEM[9970];
assign MEM[11301] = MEM[10027] + MEM[4214];
assign MEM[11302] = MEM[10031] + MEM[10016];
assign MEM[11303] = MEM[10034] + MEM[10278];
assign MEM[11304] = MEM[10036] + MEM[9883];
assign MEM[11305] = MEM[10040] + MEM[10446];
assign MEM[11306] = MEM[10043] + MEM[10238];
assign MEM[11307] = MEM[10044] + MEM[10056];
assign MEM[11308] = MEM[10048] + MEM[10181];
assign MEM[11309] = MEM[10064] + MEM[9955];
assign MEM[11310] = MEM[10093] + MEM[10321];
assign MEM[11311] = MEM[10098] + MEM[10119];
assign MEM[11312] = MEM[10103] + MEM[10113];
assign MEM[11313] = MEM[10107] + MEM[5091];
assign MEM[11314] = MEM[10111] + MEM[10136];
assign MEM[11315] = MEM[10132] + MEM[10209];
assign MEM[11316] = MEM[10146] + MEM[10193];
assign MEM[11317] = MEM[10195] + MEM[10228];
assign MEM[11318] = MEM[10198] + MEM[10012];
assign MEM[11319] = MEM[10202] + MEM[10322];
assign MEM[11320] = MEM[10205] + MEM[4731];
assign MEM[11321] = MEM[10207] + MEM[10217];
assign MEM[11322] = MEM[10218] + MEM[10112];
assign MEM[11323] = MEM[10219] + MEM[10054];
assign MEM[11324] = MEM[10269] + MEM[10192];
assign MEM[11325] = MEM[10277] + MEM[10025];
assign MEM[11326] = MEM[10408] + MEM[10286];
assign MEM[11327] = MEM[10640] + MEM[10152];
assign MEM[11328] = MEM[1415] + MEM[7359];
assign MEM[11329] = MEM[1762] + MEM[9908];
assign MEM[11330] = MEM[2327] + MEM[10167];
assign MEM[11331] = MEM[2387] + MEM[10185];
assign MEM[11332] = MEM[2805] + MEM[10150];
assign MEM[11333] = MEM[3645] + MEM[6974];
assign MEM[11334] = MEM[3687] + MEM[3698];
assign MEM[11335] = MEM[4356] + MEM[10172];
assign MEM[11336] = MEM[4533] + MEM[10079];
assign MEM[11337] = MEM[4791] + MEM[9889];
assign MEM[11338] = MEM[5067] + MEM[10389];
assign MEM[11339] = MEM[5140] + MEM[10067];
assign MEM[11340] = MEM[5493] + MEM[9943];
assign MEM[11341] = MEM[5627] + MEM[10382];
assign MEM[11342] = MEM[5684] + MEM[3349];
assign MEM[11343] = MEM[5998] + MEM[10271];
assign MEM[11344] = MEM[6291] + MEM[10397];
assign MEM[11345] = MEM[6326] + MEM[10134];
assign MEM[11346] = MEM[7239] + MEM[3519];
assign MEM[11347] = MEM[7464] + MEM[10331];
assign MEM[11348] = MEM[9676] + MEM[5426];
assign MEM[11349] = MEM[9701] + MEM[4325];
assign MEM[11350] = MEM[9736] + MEM[10024];
assign MEM[11351] = MEM[9784] + MEM[1325];
assign MEM[11352] = MEM[9825] + MEM[5671];
assign MEM[11353] = MEM[9832] + MEM[3980];
assign MEM[11354] = MEM[9879] + MEM[9915];
assign MEM[11355] = MEM[9882] + MEM[4850];
assign MEM[11356] = MEM[9919] + MEM[10039];
assign MEM[11357] = MEM[9927] + MEM[669];
assign MEM[11358] = MEM[9940] + MEM[8835];
assign MEM[11359] = MEM[9948] + MEM[3925];
assign MEM[11360] = MEM[9951] + MEM[8778];
assign MEM[11361] = MEM[9952] + MEM[2499];
assign MEM[11362] = MEM[9956] + MEM[6620];
assign MEM[11363] = MEM[9958] + MEM[6870];
assign MEM[11364] = MEM[9960] + MEM[2150];
assign MEM[11365] = MEM[9972] + MEM[1950];
assign MEM[11366] = MEM[9973] + MEM[9980];
assign MEM[11367] = MEM[9984] + MEM[5583];
assign MEM[11368] = MEM[9988] + MEM[10015];
assign MEM[11369] = MEM[9989] + MEM[10053];
assign MEM[11370] = MEM[9995] + MEM[7368];
assign MEM[11371] = MEM[10011] + MEM[4741];
assign MEM[11372] = MEM[10013] + MEM[7296];
assign MEM[11373] = MEM[10021] + MEM[4980];
assign MEM[11374] = MEM[10028] + MEM[3501];
assign MEM[11375] = MEM[10029] + MEM[4003];
assign MEM[11376] = MEM[10037] + MEM[2998];
assign MEM[11377] = MEM[10038] + MEM[3549];
assign MEM[11378] = MEM[10041] + MEM[7270];
assign MEM[11379] = MEM[10042] + MEM[3556];
assign MEM[11380] = MEM[10047] + MEM[10203];
assign MEM[11381] = MEM[10049] + MEM[3254];
assign MEM[11382] = MEM[10051] + MEM[174];
assign MEM[11383] = MEM[10060] + MEM[10155];
assign MEM[11384] = MEM[10061] + MEM[10164];
assign MEM[11385] = MEM[10063] + MEM[10080];
assign MEM[11386] = MEM[10065] + MEM[1694];
assign MEM[11387] = MEM[10066] + MEM[1341];
assign MEM[11388] = MEM[10071] + MEM[1759];
assign MEM[11389] = MEM[10072] + MEM[10086];
assign MEM[11390] = MEM[10073] + MEM[6609];
assign MEM[11391] = MEM[10074] + MEM[10105];
assign MEM[11392] = MEM[10075] + MEM[10188];
assign MEM[11393] = MEM[10076] + MEM[10114];
assign MEM[11394] = MEM[10077] + MEM[2812];
assign MEM[11395] = MEM[10078] + MEM[5246];
assign MEM[11396] = MEM[10082] + MEM[10222];
assign MEM[11397] = MEM[10085] + MEM[10307];
assign MEM[11398] = MEM[10087] + MEM[4490];
assign MEM[11399] = MEM[10088] + MEM[10233];
assign MEM[11400] = MEM[10090] + MEM[4835];
assign MEM[11401] = MEM[10092] + MEM[6180];
assign MEM[11402] = MEM[10094] + MEM[8099];
assign MEM[11403] = MEM[10095] + MEM[10169];
assign MEM[11404] = MEM[10096] + MEM[3790];
assign MEM[11405] = MEM[10100] + MEM[5910];
assign MEM[11406] = MEM[10104] + MEM[3574];
assign MEM[11407] = MEM[10106] + MEM[10006];
assign MEM[11408] = MEM[10108] + MEM[4764];
assign MEM[11409] = MEM[10110] + MEM[8219];
assign MEM[11410] = MEM[10115] + MEM[4141];
assign MEM[11411] = MEM[10116] + MEM[10214];
assign MEM[11412] = MEM[10118] + MEM[3950];
assign MEM[11413] = MEM[10120] + MEM[10186];
assign MEM[11414] = MEM[10124] + MEM[3623];
assign MEM[11415] = MEM[10126] + MEM[10206];
assign MEM[11416] = MEM[10127] + MEM[6274];
assign MEM[11417] = MEM[10129] + MEM[2510];
assign MEM[11418] = MEM[10131] + MEM[4163];
assign MEM[11419] = MEM[10133] + MEM[10316];
assign MEM[11420] = MEM[10138] + MEM[5755];
assign MEM[11421] = MEM[10141] + MEM[10176];
assign MEM[11422] = MEM[10142] + MEM[3732];
assign MEM[11423] = MEM[10143] + MEM[3302];
assign MEM[11424] = MEM[10144] + MEM[1492];
assign MEM[11425] = MEM[10145] + MEM[3447];
assign MEM[11426] = MEM[10148] + MEM[10253];
assign MEM[11427] = MEM[10153] + MEM[10161];
assign MEM[11428] = MEM[10157] + MEM[7026];
assign MEM[11429] = MEM[10158] + MEM[10480];
assign MEM[11430] = MEM[10159] + MEM[10200];
assign MEM[11431] = MEM[10160] + MEM[8212];
assign MEM[11432] = MEM[10165] + MEM[7012];
assign MEM[11433] = MEM[10166] + MEM[7619];
assign MEM[11434] = MEM[10168] + MEM[10151];
assign MEM[11435] = MEM[10170] + MEM[7498];
assign MEM[11436] = MEM[10175] + MEM[10248];
assign MEM[11437] = MEM[10184] + MEM[10215];
assign MEM[11438] = MEM[10190] + MEM[10363];
assign MEM[11439] = MEM[10191] + MEM[10208];
assign MEM[11440] = MEM[10194] + MEM[6998];
assign MEM[11441] = MEM[10196] + MEM[10287];
assign MEM[11442] = MEM[10199] + MEM[10359];
assign MEM[11443] = MEM[10204] + MEM[8636];
assign MEM[11444] = MEM[10210] + MEM[8875];
assign MEM[11445] = MEM[10211] + MEM[1076];
assign MEM[11446] = MEM[10216] + MEM[10300];
assign MEM[11447] = MEM[10224] + MEM[10282];
assign MEM[11448] = MEM[10227] + MEM[10334];
assign MEM[11449] = MEM[10229] + MEM[8742];
assign MEM[11450] = MEM[10231] + MEM[3255];
assign MEM[11451] = MEM[10234] + MEM[3003];
assign MEM[11452] = MEM[10235] + MEM[4925];
assign MEM[11453] = MEM[10236] + MEM[6170];
assign MEM[11454] = MEM[10239] + MEM[6946];
assign MEM[11455] = MEM[10240] + MEM[10427];
assign MEM[11456] = MEM[10250] + MEM[5277];
assign MEM[11457] = MEM[10252] + MEM[10350];
assign MEM[11458] = MEM[10255] + MEM[10477];
assign MEM[11459] = MEM[10256] + MEM[4254];
assign MEM[11460] = MEM[10261] + MEM[9287];
assign MEM[11461] = MEM[10263] + MEM[7394];
assign MEM[11462] = MEM[10264] + MEM[5868];
assign MEM[11463] = MEM[10268] + MEM[10365];
assign MEM[11464] = MEM[10272] + MEM[6924];
assign MEM[11465] = MEM[10273] + MEM[10242];
assign MEM[11466] = MEM[10275] + MEM[10304];
assign MEM[11467] = MEM[10276] + MEM[7283];
assign MEM[11468] = MEM[10279] + MEM[4175];
assign MEM[11469] = MEM[10288] + MEM[4589];
assign MEM[11470] = MEM[10289] + MEM[10570];
assign MEM[11471] = MEM[10295] + MEM[7762];
assign MEM[11472] = MEM[10297] + MEM[5135];
assign MEM[11473] = MEM[10298] + MEM[10342];
assign MEM[11474] = MEM[10302] + MEM[10414];
assign MEM[11475] = MEM[10306] + MEM[10459];
assign MEM[11476] = MEM[10310] + MEM[5946];
assign MEM[11477] = MEM[10315] + MEM[10246];
assign MEM[11478] = MEM[10318] + MEM[10497];
assign MEM[11479] = MEM[10319] + MEM[1254];
assign MEM[11480] = MEM[10320] + MEM[6519];
assign MEM[11481] = MEM[10326] + MEM[10343];
assign MEM[11482] = MEM[10327] + MEM[1247];
assign MEM[11483] = MEM[10332] + MEM[7603];
assign MEM[11484] = MEM[10333] + MEM[10336];
assign MEM[11485] = MEM[10337] + MEM[1172];
assign MEM[11486] = MEM[10339] + MEM[10368];
assign MEM[11487] = MEM[10341] + MEM[10571];
assign MEM[11488] = MEM[10349] + MEM[10383];
assign MEM[11489] = MEM[10353] + MEM[10424];
assign MEM[11490] = MEM[10355] + MEM[10453];
assign MEM[11491] = MEM[10357] + MEM[2946];
assign MEM[11492] = MEM[10361] + MEM[10174];
assign MEM[11493] = MEM[10366] + MEM[6286];
assign MEM[11494] = MEM[10370] + MEM[6207];
assign MEM[11495] = MEM[10376] + MEM[10464];
assign MEM[11496] = MEM[10378] + MEM[10404];
assign MEM[11497] = MEM[10381] + MEM[10399];
assign MEM[11498] = MEM[10384] + MEM[8069];
assign MEM[11499] = MEM[10385] + MEM[7260];
assign MEM[11500] = MEM[10387] + MEM[2675];
assign MEM[11501] = MEM[10391] + MEM[6271];
assign MEM[11502] = MEM[10393] + MEM[5051];
assign MEM[11503] = MEM[10395] + MEM[7101];
assign MEM[11504] = MEM[10396] + MEM[10529];
assign MEM[11505] = MEM[10402] + MEM[2165];
assign MEM[11506] = MEM[10405] + MEM[10139];
assign MEM[11507] = MEM[10407] + MEM[7847];
assign MEM[11508] = MEM[10421] + MEM[10369];
assign MEM[11509] = MEM[10430] + MEM[8836];
assign MEM[11510] = MEM[10440] + MEM[10180];
assign MEM[11511] = MEM[10452] + MEM[7590];
assign MEM[11512] = MEM[10463] + MEM[10257];
assign MEM[11513] = MEM[10498] + MEM[4359];
assign MEM[11514] = MEM[10504] + MEM[1884];
assign MEM[11515] = MEM[10515] + MEM[7428];
assign MEM[11516] = MEM[10524] + MEM[10584];
assign MEM[11517] = MEM[10526] + MEM[10827];
assign MEM[11518] = MEM[10551] + MEM[10254];
assign MEM[11519] = MEM[10558] + MEM[10266];
assign MEM[11520] = MEM[10572] + MEM[10560];
assign MEM[11521] = MEM[10594] + MEM[580];
assign MEM[11522] = MEM[10613] + MEM[1554];
assign MEM[11523] = MEM[10626] + MEM[4779];
assign MEM[11524] = MEM[10666] + MEM[2395];
assign MEM[11525] = MEM[10684] + MEM[1813];
assign MEM[11526] = MEM[10701] + MEM[1367];
assign MEM[11527] = MEM[101] + MEM[7928];
assign MEM[11528] = MEM[135] + MEM[10371];
assign MEM[11529] = MEM[230] + MEM[5107];
assign MEM[11530] = MEM[263] + MEM[2101];
assign MEM[11531] = MEM[276] + MEM[10232];
assign MEM[11532] = MEM[286] + MEM[10512];
assign MEM[11533] = MEM[357] + MEM[10293];
assign MEM[11534] = MEM[370] + MEM[830];
assign MEM[11535] = MEM[372] + MEM[10329];
assign MEM[11536] = MEM[399] + MEM[1015];
assign MEM[11537] = MEM[414] + MEM[1094];
assign MEM[11538] = MEM[423] + MEM[10587];
assign MEM[11539] = MEM[479] + MEM[10348];
assign MEM[11540] = MEM[503] + MEM[10344];
assign MEM[11541] = MEM[519] + MEM[9055];
assign MEM[11542] = MEM[522] + MEM[10084];
assign MEM[11543] = MEM[524] + MEM[5231];
assign MEM[11544] = MEM[549] + MEM[7658];
assign MEM[11545] = MEM[589] + MEM[10283];
assign MEM[11546] = MEM[610] + MEM[8060];
assign MEM[11547] = MEM[635] + MEM[4542];
assign MEM[11548] = MEM[647] + MEM[10367];
assign MEM[11549] = MEM[710] + MEM[1548];
assign MEM[11550] = MEM[746] + MEM[3845];
assign MEM[11551] = MEM[770] + MEM[5527];
assign MEM[11552] = MEM[781] + MEM[6109];
assign MEM[11553] = MEM[790] + MEM[10372];
assign MEM[11554] = MEM[795] + MEM[10501];
assign MEM[11555] = MEM[806] + MEM[8669];
assign MEM[11556] = MEM[813] + MEM[10284];
assign MEM[11557] = MEM[822] + MEM[10323];
assign MEM[11558] = MEM[823] + MEM[1301];
assign MEM[11559] = MEM[942] + MEM[10443];
assign MEM[11560] = MEM[956] + MEM[7729];
assign MEM[11561] = MEM[989] + MEM[1708];
assign MEM[11562] = MEM[1023] + MEM[1772];
assign MEM[11563] = MEM[1044] + MEM[8607];
assign MEM[11564] = MEM[1046] + MEM[7217];
assign MEM[11565] = MEM[1054] + MEM[5420];
assign MEM[11566] = MEM[1084] + MEM[2918];
assign MEM[11567] = MEM[1125] + MEM[2700];
assign MEM[11568] = MEM[1173] + MEM[10265];
assign MEM[11569] = MEM[1181] + MEM[5323];
assign MEM[11570] = MEM[1238] + MEM[10156];
assign MEM[11571] = MEM[1262] + MEM[6681];
assign MEM[11572] = MEM[1293] + MEM[7851];
assign MEM[11573] = MEM[1358] + MEM[2207];
assign MEM[11574] = MEM[1363] + MEM[2836];
assign MEM[11575] = MEM[1364] + MEM[10696];
assign MEM[11576] = MEM[1403] + MEM[2461];
assign MEM[11577] = MEM[1412] + MEM[7719];
assign MEM[11578] = MEM[1426] + MEM[8108];
assign MEM[11579] = MEM[1447] + MEM[10154];
assign MEM[11580] = MEM[1470] + MEM[1303];
assign MEM[11581] = MEM[1475] + MEM[6913];
assign MEM[11582] = MEM[1502] + MEM[9614];
assign MEM[11583] = MEM[1518] + MEM[5541];
assign MEM[11584] = MEM[1575] + MEM[10468];
assign MEM[11585] = MEM[1581] + MEM[10410];
assign MEM[11586] = MEM[1591] + MEM[10400];
assign MEM[11587] = MEM[1717] + MEM[10589];
assign MEM[11588] = MEM[1719] + MEM[2571];
assign MEM[11589] = MEM[1763] + MEM[2685];
assign MEM[11590] = MEM[1788] + MEM[5459];
assign MEM[11591] = MEM[1805] + MEM[3691];
assign MEM[11592] = MEM[1820] + MEM[4390];
assign MEM[11593] = MEM[1826] + MEM[10451];
assign MEM[11594] = MEM[1835] + MEM[4588];
assign MEM[11595] = MEM[1886] + MEM[10220];
assign MEM[11596] = MEM[1914] + MEM[10375];
assign MEM[11597] = MEM[1947] + MEM[1782];
assign MEM[11598] = MEM[1948] + MEM[7102];
assign MEM[11599] = MEM[2004] + MEM[5754];
assign MEM[11600] = MEM[2011] + MEM[5914];
assign MEM[11601] = MEM[2030] + MEM[10294];
assign MEM[11602] = MEM[2063] + MEM[3603];
assign MEM[11603] = MEM[2079] + MEM[7268];
assign MEM[11604] = MEM[2082] + MEM[5708];
assign MEM[11605] = MEM[2123] + MEM[5907];
assign MEM[11606] = MEM[2171] + MEM[10555];
assign MEM[11607] = MEM[2175] + MEM[10099];
assign MEM[11608] = MEM[2198] + MEM[7162];
assign MEM[11609] = MEM[2210] + MEM[2716];
assign MEM[11610] = MEM[2282] + MEM[8653];
assign MEM[11611] = MEM[2293] + MEM[6385];
assign MEM[11612] = MEM[2326] + MEM[10447];
assign MEM[11613] = MEM[2340] + MEM[6038];
assign MEM[11614] = MEM[2397] + MEM[2766];
assign MEM[11615] = MEM[2423] + MEM[10521];
assign MEM[11616] = MEM[2427] + MEM[5815];
assign MEM[11617] = MEM[2431] + MEM[6967];
assign MEM[11618] = MEM[2470] + MEM[10476];
assign MEM[11619] = MEM[2500] + MEM[3661];
assign MEM[11620] = MEM[2535] + MEM[10358];
assign MEM[11621] = MEM[2613] + MEM[8654];
assign MEM[11622] = MEM[2652] + MEM[10409];
assign MEM[11623] = MEM[2748] + MEM[10178];
assign MEM[11624] = MEM[2759] + MEM[5863];
assign MEM[11625] = MEM[2838] + MEM[10345];
assign MEM[11626] = MEM[2859] + MEM[3679];
assign MEM[11627] = MEM[2866] + MEM[3422];
assign MEM[11628] = MEM[2871] + MEM[6685];
assign MEM[11629] = MEM[2894] + MEM[5027];
assign MEM[11630] = MEM[2899] + MEM[10422];
assign MEM[11631] = MEM[2910] + MEM[6119];
assign MEM[11632] = MEM[2954] + MEM[5727];
assign MEM[11633] = MEM[2987] + MEM[10171];
assign MEM[11634] = MEM[3029] + MEM[10230];
assign MEM[11635] = MEM[3047] + MEM[2235];
assign MEM[11636] = MEM[3067] + MEM[10325];
assign MEM[11637] = MEM[3087] + MEM[9398];
assign MEM[11638] = MEM[3091] + MEM[10455];
assign MEM[11639] = MEM[3125] + MEM[10482];
assign MEM[11640] = MEM[3167] + MEM[10259];
assign MEM[11641] = MEM[3182] + MEM[7784];
assign MEM[11642] = MEM[3220] + MEM[10628];
assign MEM[11643] = MEM[3228] + MEM[6822];
assign MEM[11644] = MEM[3247] + MEM[4941];
assign MEM[11645] = MEM[3250] + MEM[10392];
assign MEM[11646] = MEM[3311] + MEM[6915];
assign MEM[11647] = MEM[3327] + MEM[10281];
assign MEM[11648] = MEM[3346] + MEM[6996];
assign MEM[11649] = MEM[3347] + MEM[7246];
assign MEM[11650] = MEM[3386] + MEM[10135];
assign MEM[11651] = MEM[3389] + MEM[10121];
assign MEM[11652] = MEM[3399] + MEM[2386];
assign MEM[11653] = MEM[3420] + MEM[8411];
assign MEM[11654] = MEM[3439] + MEM[10563];
assign MEM[11655] = MEM[3468] + MEM[6429];
assign MEM[11656] = MEM[3491] + MEM[10362];
assign MEM[11657] = MEM[3493] + MEM[10496];
assign MEM[11658] = MEM[3651] + MEM[1090];
assign MEM[11659] = MEM[3662] + MEM[5311];
assign MEM[11660] = MEM[3671] + MEM[10522];
assign MEM[11661] = MEM[3675] + MEM[10221];
assign MEM[11662] = MEM[3684] + MEM[9000];
assign MEM[11663] = MEM[3701] + MEM[10454];
assign MEM[11664] = MEM[3719] + MEM[6966];
assign MEM[11665] = MEM[3724] + MEM[11021];
assign MEM[11666] = MEM[3754] + MEM[6493];
assign MEM[11667] = MEM[3765] + MEM[1828];
assign MEM[11668] = MEM[3855] + MEM[6741];
assign MEM[11669] = MEM[3894] + MEM[2994];
assign MEM[11670] = MEM[3927] + MEM[7388];
assign MEM[11671] = MEM[3957] + MEM[4066];
assign MEM[11672] = MEM[3963] + MEM[3743];
assign MEM[11673] = MEM[3967] + MEM[3141];
assign MEM[11674] = MEM[3987] + MEM[3839];
assign MEM[11675] = MEM[4030] + MEM[6683];
assign MEM[11676] = MEM[4038] + MEM[6518];
assign MEM[11677] = MEM[4068] + MEM[6127];
assign MEM[11678] = MEM[4094] + MEM[573];
assign MEM[11679] = MEM[4103] + MEM[10290];
assign MEM[11680] = MEM[4130] + MEM[5333];
assign MEM[11681] = MEM[4167] + MEM[10243];
assign MEM[11682] = MEM[4190] + MEM[845];
assign MEM[11683] = MEM[4219] + MEM[10516];
assign MEM[11684] = MEM[4226] + MEM[10426];
assign MEM[11685] = MEM[4262] + MEM[4951];
assign MEM[11686] = MEM[4263] + MEM[2837];
assign MEM[11687] = MEM[4294] + MEM[5621];
assign MEM[11688] = MEM[4342] + MEM[4668];
assign MEM[11689] = MEM[4350] + MEM[10356];
assign MEM[11690] = MEM[4351] + MEM[2821];
assign MEM[11691] = MEM[4366] + MEM[8641];
assign MEM[11692] = MEM[4374] + MEM[10225];
assign MEM[11693] = MEM[4389] + MEM[6378];
assign MEM[11694] = MEM[4414] + MEM[4667];
assign MEM[11695] = MEM[4419] + MEM[9632];
assign MEM[11696] = MEM[4455] + MEM[10237];
assign MEM[11697] = MEM[4461] + MEM[9019];
assign MEM[11698] = MEM[4510] + MEM[5933];
assign MEM[11699] = MEM[4578] + MEM[10491];
assign MEM[11700] = MEM[4596] + MEM[2607];
assign MEM[11701] = MEM[4606] + MEM[8371];
assign MEM[11702] = MEM[4629] + MEM[9396];
assign MEM[11703] = MEM[4630] + MEM[3903];
assign MEM[11704] = MEM[4635] + MEM[2562];
assign MEM[11705] = MEM[4659] + MEM[5973];
assign MEM[11706] = MEM[4660] + MEM[3083];
assign MEM[11707] = MEM[4687] + MEM[215];
assign MEM[11708] = MEM[4693] + MEM[5996];
assign MEM[11709] = MEM[4703] + MEM[10373];
assign MEM[11710] = MEM[4732] + MEM[8395];
assign MEM[11711] = MEM[4734] + MEM[10434];
assign MEM[11712] = MEM[4746] + MEM[6863];
assign MEM[11713] = MEM[4804] + MEM[10532];
assign MEM[11714] = MEM[4807] + MEM[10401];
assign MEM[11715] = MEM[4815] + MEM[6806];
assign MEM[11716] = MEM[4831] + MEM[10244];
assign MEM[11717] = MEM[4837] + MEM[8206];
assign MEM[11718] = MEM[4842] + MEM[941];
assign MEM[11719] = MEM[4878] + MEM[2786];
assign MEM[11720] = MEM[4891] + MEM[494];
assign MEM[11721] = MEM[4943] + MEM[10352];
assign MEM[11722] = MEM[4957] + MEM[10296];
assign MEM[11723] = MEM[4991] + MEM[10542];
assign MEM[11724] = MEM[4995] + MEM[10543];
assign MEM[11725] = MEM[5031] + MEM[10456];
assign MEM[11726] = MEM[5095] + MEM[6022];
assign MEM[11727] = MEM[5122] + MEM[3286];
assign MEM[11728] = MEM[5150] + MEM[7979];
assign MEM[11729] = MEM[5165] + MEM[7811];
assign MEM[11730] = MEM[5171] + MEM[8433];
assign MEM[11731] = MEM[5175] + MEM[4316];
assign MEM[11732] = MEM[5238] + MEM[5725];
assign MEM[11733] = MEM[5247] + MEM[2419];
assign MEM[11734] = MEM[5268] + MEM[125];
assign MEM[11735] = MEM[5293] + MEM[10245];
assign MEM[11736] = MEM[5306] + MEM[6283];
assign MEM[11737] = MEM[5307] + MEM[1999];
assign MEM[11738] = MEM[5308] + MEM[10262];
assign MEM[11739] = MEM[5310] + MEM[8011];
assign MEM[11740] = MEM[5317] + MEM[1446];
assign MEM[11741] = MEM[5354] + MEM[4031];
assign MEM[11742] = MEM[5358] + MEM[3423];
assign MEM[11743] = MEM[5365] + MEM[10258];
assign MEM[11744] = MEM[5373] + MEM[2839];
assign MEM[11745] = MEM[5374] + MEM[10137];
assign MEM[11746] = MEM[5389] + MEM[7133];
assign MEM[11747] = MEM[5396] + MEM[3276];
assign MEM[11748] = MEM[5398] + MEM[4275];
assign MEM[11749] = MEM[5412] + MEM[6423];
assign MEM[11750] = MEM[5414] + MEM[3750];
assign MEM[11751] = MEM[5437] + MEM[10417];
assign MEM[11752] = MEM[5485] + MEM[7382];
assign MEM[11753] = MEM[5518] + MEM[7407];
assign MEM[11754] = MEM[5535] + MEM[4100];
assign MEM[11755] = MEM[5548] + MEM[10420];
assign MEM[11756] = MEM[5557] + MEM[5559];
assign MEM[11757] = MEM[5597] + MEM[5510];
assign MEM[11758] = MEM[5614] + MEM[1892];
assign MEM[11759] = MEM[5668] + MEM[1213];
assign MEM[11760] = MEM[5701] + MEM[1660];
assign MEM[11761] = MEM[5716] + MEM[6002];
assign MEM[11762] = MEM[5719] + MEM[2942];
assign MEM[11763] = MEM[5724] + MEM[8222];
assign MEM[11764] = MEM[5730] + MEM[10189];
assign MEM[11765] = MEM[5796] + MEM[6975];
assign MEM[11766] = MEM[5799] + MEM[2883];
assign MEM[11767] = MEM[5822] + MEM[8479];
assign MEM[11768] = MEM[5854] + MEM[5901];
assign MEM[11769] = MEM[5875] + MEM[4286];
assign MEM[11770] = MEM[5882] + MEM[5251];
assign MEM[11771] = MEM[5926] + MEM[7626];
assign MEM[11772] = MEM[5927] + MEM[3437];
assign MEM[11773] = MEM[5936] + MEM[2875];
assign MEM[11774] = MEM[5949] + MEM[7922];
assign MEM[11775] = MEM[5955] + MEM[7216];
assign MEM[11776] = MEM[5957] + MEM[7930];
assign MEM[11777] = MEM[5963] + MEM[1778];
assign MEM[11778] = MEM[5978] + MEM[10518];
assign MEM[11779] = MEM[5987] + MEM[10442];
assign MEM[11780] = MEM[5999] + MEM[7528];
assign MEM[11781] = MEM[6006] + MEM[10416];
assign MEM[11782] = MEM[6014] + MEM[2071];
assign MEM[11783] = MEM[6063] + MEM[5958];
assign MEM[11784] = MEM[6070] + MEM[10441];
assign MEM[11785] = MEM[6077] + MEM[6436];
assign MEM[11786] = MEM[6095] + MEM[2959];
assign MEM[11787] = MEM[6118] + MEM[5103];
assign MEM[11788] = MEM[6130] + MEM[287];
assign MEM[11789] = MEM[6149] + MEM[10314];
assign MEM[11790] = MEM[6151] + MEM[2074];
assign MEM[11791] = MEM[6183] + MEM[10299];
assign MEM[11792] = MEM[6197] + MEM[6515];
assign MEM[11793] = MEM[6273] + MEM[10374];
assign MEM[11794] = MEM[6288] + MEM[2277];
assign MEM[11795] = MEM[6295] + MEM[5573];
assign MEM[11796] = MEM[6296] + MEM[10102];
assign MEM[11797] = MEM[6300] + MEM[7520];
assign MEM[11798] = MEM[6301] + MEM[5791];
assign MEM[11799] = MEM[6310] + MEM[10364];
assign MEM[11800] = MEM[6315] + MEM[4117];
assign MEM[11801] = MEM[6327] + MEM[8315];
assign MEM[11802] = MEM[6418] + MEM[10241];
assign MEM[11803] = MEM[6427] + MEM[8144];
assign MEM[11804] = MEM[6441] + MEM[4199];
assign MEM[11805] = MEM[6446] + MEM[2355];
assign MEM[11806] = MEM[6467] + MEM[5599];
assign MEM[11807] = MEM[6468] + MEM[7086];
assign MEM[11808] = MEM[6471] + MEM[555];
assign MEM[11809] = MEM[6561] + MEM[7577];
assign MEM[11810] = MEM[6658] + MEM[10415];
assign MEM[11811] = MEM[6693] + MEM[3133];
assign MEM[11812] = MEM[6710] + MEM[6279];
assign MEM[11813] = MEM[6718] + MEM[1029];
assign MEM[11814] = MEM[6774] + MEM[3306];
assign MEM[11815] = MEM[6797] + MEM[603];
assign MEM[11816] = MEM[6803] + MEM[7685];
assign MEM[11817] = MEM[6810] + MEM[6230];
assign MEM[11818] = MEM[6826] + MEM[2930];
assign MEM[11819] = MEM[6832] + MEM[8816];
assign MEM[11820] = MEM[6856] + MEM[10338];
assign MEM[11821] = MEM[6876] + MEM[7305];
assign MEM[11822] = MEM[6908] + MEM[6776];
assign MEM[11823] = MEM[6954] + MEM[9693];
assign MEM[11824] = MEM[6962] + MEM[10301];
assign MEM[11825] = MEM[6976] + MEM[10460];
assign MEM[11826] = MEM[7013] + MEM[8111];
assign MEM[11827] = MEM[7019] + MEM[6223];
assign MEM[11828] = MEM[7028] + MEM[6299];
assign MEM[11829] = MEM[7029] + MEM[10535];
assign MEM[11830] = MEM[7051] + MEM[902];
assign MEM[11831] = MEM[7053] + MEM[7126];
assign MEM[11832] = MEM[7073] + MEM[6037];
assign MEM[11833] = MEM[7108] + MEM[10583];
assign MEM[11834] = MEM[7129] + MEM[7573];
assign MEM[11835] = MEM[7130] + MEM[7234];
assign MEM[11836] = MEM[7140] + MEM[10514];
assign MEM[11837] = MEM[7178] + MEM[9792];
assign MEM[11838] = MEM[7207] + MEM[10562];
assign MEM[11839] = MEM[7209] + MEM[4020];
assign MEM[11840] = MEM[7252] + MEM[8146];
assign MEM[11841] = MEM[7272] + MEM[1932];
assign MEM[11842] = MEM[7299] + MEM[10097];
assign MEM[11843] = MEM[7380] + MEM[8890];
assign MEM[11844] = MEM[7624] + MEM[10568];
assign MEM[11845] = MEM[7627] + MEM[8347];
assign MEM[11846] = MEM[7650] + MEM[6386];
assign MEM[11847] = MEM[7693] + MEM[10634];
assign MEM[11848] = MEM[7722] + MEM[10285];
assign MEM[11849] = MEM[7736] + MEM[1695];
assign MEM[11850] = MEM[7780] + MEM[4909];
assign MEM[11851] = MEM[7805] + MEM[8119];
assign MEM[11852] = MEM[7819] + MEM[10490];
assign MEM[11853] = MEM[7899] + MEM[4004];
assign MEM[11854] = MEM[7924] + MEM[10412];
assign MEM[11855] = MEM[7960] + MEM[2269];
assign MEM[11856] = MEM[8058] + MEM[5971];
assign MEM[11857] = MEM[8089] + MEM[10212];
assign MEM[11858] = MEM[8123] + MEM[10386];
assign MEM[11859] = MEM[8295] + MEM[10303];
assign MEM[11860] = MEM[8333] + MEM[1775];
assign MEM[11861] = MEM[8488] + MEM[8929];
assign MEM[11862] = MEM[8551] + MEM[6928];
assign MEM[11863] = MEM[8676] + MEM[7778];
assign MEM[11864] = MEM[8805] + MEM[10707];
assign MEM[11865] = MEM[8886] + MEM[7039];
assign MEM[11866] = MEM[8995] + MEM[8790];
assign MEM[11867] = MEM[9178] + MEM[9754];
assign MEM[11868] = MEM[9241] + MEM[9430];
assign MEM[11869] = MEM[9275] + MEM[10680];
assign MEM[11870] = MEM[9454] + MEM[10470];
assign MEM[11871] = MEM[9458] + MEM[1946];
assign MEM[11872] = MEM[9486] + MEM[4447];
assign MEM[11873] = MEM[9653] + MEM[1797];
assign MEM[11874] = MEM[9860] + MEM[10679];
assign MEM[11875] = MEM[10062] + MEM[317];
assign MEM[11876] = MEM[10081] + MEM[1750];
assign MEM[11877] = MEM[10091] + MEM[2159];
assign MEM[11878] = MEM[10182] + MEM[2084];
assign MEM[11879] = MEM[10183] + MEM[670];
assign MEM[11880] = MEM[10223] + MEM[6909];
assign MEM[11881] = MEM[10226] + MEM[3469];
assign MEM[11882] = MEM[10249] + MEM[2667];
assign MEM[11883] = MEM[10251] + MEM[10457];
assign MEM[11884] = MEM[10260] + MEM[7370];
assign MEM[11885] = MEM[10267] + MEM[3078];
assign MEM[11886] = MEM[10270] + MEM[6582];
assign MEM[11887] = MEM[10274] + MEM[254];
assign MEM[11888] = MEM[10280] + MEM[5678];
assign MEM[11889] = MEM[10291] + MEM[971];
assign MEM[11890] = MEM[10305] + MEM[3542];
assign MEM[11891] = MEM[10308] + MEM[7257];
assign MEM[11892] = MEM[10309] + MEM[3495];
assign MEM[11893] = MEM[10311] + MEM[6705];
assign MEM[11894] = MEM[10312] + MEM[3902];
assign MEM[11895] = MEM[10313] + MEM[1252];
assign MEM[11896] = MEM[10317] + MEM[1093];
assign MEM[11897] = MEM[10324] + MEM[5173];
assign MEM[11898] = MEM[10328] + MEM[2258];
assign MEM[11899] = MEM[10335] + MEM[4565];
assign MEM[11900] = MEM[10340] + MEM[725];
assign MEM[11901] = MEM[10346] + MEM[5531];
assign MEM[11902] = MEM[10347] + MEM[4701];
assign MEM[11903] = MEM[10351] + MEM[4655];
assign MEM[11904] = MEM[10354] + MEM[2982];
assign MEM[11905] = MEM[10360] + MEM[30];
assign MEM[11906] = MEM[10377] + MEM[775];
assign MEM[11907] = MEM[10380] + MEM[4607];
assign MEM[11908] = MEM[10388] + MEM[1270];
assign MEM[11909] = MEM[10390] + MEM[10481];
assign MEM[11910] = MEM[10394] + MEM[4573];
assign MEM[11911] = MEM[10398] + MEM[3517];
assign MEM[11912] = MEM[10403] + MEM[3429];
assign MEM[11913] = MEM[10406] + MEM[1189];
assign MEM[11914] = MEM[10411] + MEM[7201];
assign MEM[11915] = MEM[10413] + MEM[10520];
assign MEM[11916] = MEM[10418] + MEM[2206];
assign MEM[11917] = MEM[10419] + MEM[581];
assign MEM[11918] = MEM[10423] + MEM[5925];
assign MEM[11919] = MEM[10425] + MEM[10552];
assign MEM[11920] = MEM[10428] + MEM[7857];
assign MEM[11921] = MEM[10429] + MEM[10629];
assign MEM[11922] = MEM[10431] + MEM[10511];
assign MEM[11923] = MEM[10432] + MEM[2428];
assign MEM[11924] = MEM[10433] + MEM[3983];
assign MEM[11925] = MEM[10435] + MEM[5539];
assign MEM[11926] = MEM[10436] + MEM[1677];
assign MEM[11927] = MEM[10438] + MEM[4718];
assign MEM[11928] = MEM[10439] + MEM[5074];
assign MEM[11929] = MEM[10444] + MEM[3367];
assign MEM[11930] = MEM[10448] + MEM[548];
assign MEM[11931] = MEM[10449] + MEM[2444];
assign MEM[11932] = MEM[10450] + MEM[5487];
assign MEM[11933] = MEM[10458] + MEM[10510];
assign MEM[11934] = MEM[10461] + MEM[4987];
assign MEM[11935] = MEM[10465] + MEM[2451];
assign MEM[11936] = MEM[10467] + MEM[7273];
assign MEM[11937] = MEM[10469] + MEM[7116];
assign MEM[11938] = MEM[10471] + MEM[6175];
assign MEM[11939] = MEM[10472] + MEM[3085];
assign MEM[11940] = MEM[10473] + MEM[1157];
assign MEM[11941] = MEM[10474] + MEM[118];
assign MEM[11942] = MEM[10475] + MEM[3340];
assign MEM[11943] = MEM[10478] + MEM[4964];
assign MEM[11944] = MEM[10479] + MEM[3676];
assign MEM[11945] = MEM[10483] + MEM[2715];
assign MEM[11946] = MEM[10484] + MEM[10528];
assign MEM[11947] = MEM[10485] + MEM[7238];
assign MEM[11948] = MEM[10486] + MEM[2605];
assign MEM[11949] = MEM[10488] + MEM[5853];
assign MEM[11950] = MEM[10489] + MEM[141];
assign MEM[11951] = MEM[10492] + MEM[5055];
assign MEM[11952] = MEM[10493] + MEM[2438];
assign MEM[11953] = MEM[10494] + MEM[6062];
assign MEM[11954] = MEM[10495] + MEM[3565];
assign MEM[11955] = MEM[10499] + MEM[10567];
assign MEM[11956] = MEM[10502] + MEM[1770];
assign MEM[11957] = MEM[10503] + MEM[151];
assign MEM[11958] = MEM[10505] + MEM[10668];
assign MEM[11959] = MEM[10506] + MEM[10599];
assign MEM[11960] = MEM[10507] + MEM[2917];
assign MEM[11961] = MEM[10508] + MEM[10610];
assign MEM[11962] = MEM[10509] + MEM[3981];
assign MEM[11963] = MEM[10513] + MEM[10527];
assign MEM[11964] = MEM[10517] + MEM[10561];
assign MEM[11965] = MEM[10519] + MEM[3653];
assign MEM[11966] = MEM[10523] + MEM[8743];
assign MEM[11967] = MEM[10525] + MEM[4444];
assign MEM[11968] = MEM[10533] + MEM[2924];
assign MEM[11969] = MEM[10534] + MEM[8887];
assign MEM[11970] = MEM[10536] + MEM[10553];
assign MEM[11971] = MEM[10537] + MEM[7943];
assign MEM[11972] = MEM[10538] + MEM[333];
assign MEM[11973] = MEM[10539] + MEM[245];
assign MEM[11974] = MEM[10540] + MEM[8830];
assign MEM[11975] = MEM[10541] + MEM[523];
assign MEM[11976] = MEM[10544] + MEM[541];
assign MEM[11977] = MEM[10546] + MEM[2574];
assign MEM[11978] = MEM[10547] + MEM[2901];
assign MEM[11979] = MEM[10548] + MEM[4695];
assign MEM[11980] = MEM[10549] + MEM[6804];
assign MEM[11981] = MEM[10550] + MEM[6229];
assign MEM[11982] = MEM[10554] + MEM[3829];
assign MEM[11983] = MEM[10556] + MEM[7403];
assign MEM[11984] = MEM[10557] + MEM[10611];
assign MEM[11985] = MEM[10564] + MEM[1930];
assign MEM[11986] = MEM[10566] + MEM[8746];
assign MEM[11987] = MEM[10579] + MEM[2180];
assign MEM[11988] = MEM[10588] + MEM[8217];
assign MEM[11989] = MEM[10592] + MEM[1860];
assign MEM[11990] = MEM[10596] + MEM[2546];
assign MEM[11991] = MEM[10597] + MEM[3866];
assign MEM[11992] = MEM[10601] + MEM[2077];
assign MEM[11993] = MEM[10604] + MEM[731];
assign MEM[11994] = MEM[10614] + MEM[355];
assign MEM[11995] = MEM[10617] + MEM[8311];
assign MEM[11996] = MEM[10618] + MEM[4739];
assign MEM[11997] = MEM[10620] + MEM[6579];
assign MEM[11998] = MEM[10622] + MEM[8775];
assign MEM[11999] = MEM[10625] + MEM[1654];
assign MEM[12000] = MEM[10630] + MEM[10643];
assign MEM[12001] = MEM[10632] + MEM[3031];
assign MEM[12002] = MEM[10636] + MEM[5924];
assign MEM[12003] = MEM[10637] + MEM[351];
assign MEM[12004] = MEM[10641] + MEM[5471];
assign MEM[12005] = MEM[10646] + MEM[1004];
assign MEM[12006] = MEM[10647] + MEM[3551];
assign MEM[12007] = MEM[10648] + MEM[3099];
assign MEM[12008] = MEM[10650] + MEM[556];
assign MEM[12009] = MEM[10651] + MEM[8569];
assign MEM[12010] = MEM[10652] + MEM[955];
assign MEM[12011] = MEM[10653] + MEM[8915];
assign MEM[12012] = MEM[10654] + MEM[3463];
assign MEM[12013] = MEM[10657] + MEM[366];
assign MEM[12014] = MEM[10661] + MEM[6078];
assign MEM[12015] = MEM[10662] + MEM[7835];
assign MEM[12016] = MEM[10663] + MEM[1821];
assign MEM[12017] = MEM[10665] + MEM[7800];
assign MEM[12018] = MEM[10669] + MEM[3990];
assign MEM[12019] = MEM[10670] + MEM[255];
assign MEM[12020] = MEM[10673] + MEM[6667];
assign MEM[12021] = MEM[10676] + MEM[405];
assign MEM[12022] = MEM[10677] + MEM[3835];
assign MEM[12023] = MEM[10683] + MEM[5756];
assign MEM[12024] = MEM[10686] + MEM[3834];
assign MEM[12025] = MEM[10687] + MEM[4519];
assign MEM[12026] = MEM[10689] + MEM[901];
assign MEM[12027] = MEM[10690] + MEM[4853];
assign MEM[12028] = MEM[10695] + MEM[6470];
assign MEM[12029] = MEM[10698] + MEM[643];
assign MEM[12030] = MEM[10700] + MEM[516];
assign MEM[12031] = MEM[10702] + MEM[1798];
assign MEM[12032] = MEM[10703] + MEM[3357];
assign MEM[12033] = MEM[10704] + MEM[5909];
assign MEM[12034] = MEM[10706] + MEM[10761];
assign MEM[12035] = MEM[10709] + MEM[8576];
assign MEM[12036] = MEM[10711] + MEM[4197];
assign MEM[12037] = MEM[10713] + MEM[2477];
assign MEM[12038] = MEM[10719] + MEM[5846];
assign MEM[12039] = MEM[10722] + MEM[2734];
assign MEM[12040] = MEM[10729] + MEM[10789];
assign MEM[12041] = MEM[10731] + MEM[6565];
assign MEM[12042] = MEM[10732] + MEM[8606];
assign MEM[12043] = MEM[10734] + MEM[10795];
assign MEM[12044] = MEM[10736] + MEM[3479];
assign MEM[12045] = MEM[10740] + MEM[3582];
assign MEM[12046] = MEM[10764] + MEM[1428];
assign MEM[12047] = MEM[10766] + MEM[11117];
assign MEM[12048] = MEM[10767] + MEM[7598];
assign MEM[12049] = MEM[10777] + MEM[6372];
assign MEM[12050] = MEM[10794] + MEM[8057];
assign MEM[12051] = MEM[10799] + MEM[4210];
assign MEM[12052] = MEM[10813] + MEM[5204];
assign MEM[12053] = MEM[10824] + MEM[1731];
assign MEM[12054] = MEM[10832] + MEM[5580];
assign MEM[12055] = MEM[10835] + MEM[1606];
assign MEM[12056] = MEM[10839] + MEM[7020];
assign MEM[12057] = MEM[10849] + MEM[10741];
assign MEM[12058] = MEM[10850] + MEM[308];
assign MEM[12059] = MEM[10864] + MEM[4339];
assign MEM[12060] = MEM[10865] + MEM[818];
assign MEM[12061] = MEM[10874] + MEM[6289];
assign MEM[12062] = MEM[10877] + MEM[3023];
assign MEM[12063] = MEM[10878] + MEM[7059];
assign MEM[12064] = MEM[10883] + MEM[2902];
assign MEM[12065] = MEM[10924] + MEM[5108];
assign MEM[12066] = MEM[10927] + MEM[4147];
assign MEM[12067] = MEM[10941] + MEM[3214];
assign MEM[12068] = MEM[10954] + MEM[10655];
assign MEM[12069] = MEM[10960] + MEM[8258];
assign MEM[12070] = MEM[10995] + MEM[8231];
assign MEM[12071] = MEM[11008] + MEM[5661];
assign MEM[12072] = MEM[11019] + MEM[6617];
assign MEM[12073] = MEM[5] + MEM[7046];
assign MEM[12074] = MEM[6] + MEM[4557];
assign MEM[12075] = MEM[13] + MEM[5943];
assign MEM[12076] = MEM[14] + MEM[4013];
assign MEM[12077] = MEM[15] + MEM[6444];
assign MEM[12078] = MEM[21] + MEM[3101];
assign MEM[12079] = MEM[22] + MEM[6945];
assign MEM[12080] = MEM[23] + MEM[2541];
assign MEM[12081] = MEM[29] + MEM[2109];
assign MEM[12082] = MEM[37] + MEM[2669];
assign MEM[12083] = MEM[39] + MEM[10615];
assign MEM[12084] = MEM[45] + MEM[614];
assign MEM[12085] = MEM[46] + MEM[526];
assign MEM[12086] = MEM[70] + MEM[1823];
assign MEM[12087] = MEM[77] + MEM[6311];
assign MEM[12088] = MEM[86] + MEM[2981];
assign MEM[12089] = MEM[87] + MEM[5607];
assign MEM[12090] = MEM[95] + MEM[4253];
assign MEM[12091] = MEM[117] + MEM[7500];
assign MEM[12092] = MEM[126] + MEM[7249];
assign MEM[12093] = MEM[127] + MEM[3780];
assign MEM[12094] = MEM[134] + MEM[5267];
assign MEM[12095] = MEM[149] + MEM[5054];
assign MEM[12096] = MEM[159] + MEM[1487];
assign MEM[12097] = MEM[165] + MEM[5356];
assign MEM[12098] = MEM[175] + MEM[3309];
assign MEM[12099] = MEM[183] + MEM[970];
assign MEM[12100] = MEM[189] + MEM[6477];
assign MEM[12101] = MEM[190] + MEM[1644];
assign MEM[12102] = MEM[198] + MEM[10437];
assign MEM[12103] = MEM[199] + MEM[2299];
assign MEM[12104] = MEM[207] + MEM[2661];
assign MEM[12105] = MEM[221] + MEM[1519];
assign MEM[12106] = MEM[222] + MEM[7687];
assign MEM[12107] = MEM[231] + MEM[9155];
assign MEM[12108] = MEM[237] + MEM[269];
assign MEM[12109] = MEM[239] + MEM[1020];
assign MEM[12110] = MEM[247] + MEM[7750];
assign MEM[12111] = MEM[271] + MEM[1237];
assign MEM[12112] = MEM[277] + MEM[2637];
assign MEM[12113] = MEM[279] + MEM[1290];
assign MEM[12114] = MEM[284] + MEM[915];
assign MEM[12115] = MEM[293] + MEM[870];
assign MEM[12116] = MEM[294] + MEM[4562];
assign MEM[12117] = MEM[295] + MEM[991];
assign MEM[12118] = MEM[301] + MEM[5438];
assign MEM[12119] = MEM[302] + MEM[3293];
assign MEM[12120] = MEM[307] + MEM[1243];
assign MEM[12121] = MEM[309] + MEM[1963];
assign MEM[12122] = MEM[310] + MEM[9765];
assign MEM[12123] = MEM[311] + MEM[7532];
assign MEM[12124] = MEM[315] + MEM[1087];
assign MEM[12125] = MEM[316] + MEM[756];
assign MEM[12126] = MEM[318] + MEM[4442];
assign MEM[12127] = MEM[323] + MEM[2723];
assign MEM[12128] = MEM[324] + MEM[1431];
assign MEM[12129] = MEM[330] + MEM[4306];
assign MEM[12130] = MEM[332] + MEM[1924];
assign MEM[12131] = MEM[334] + MEM[2092];
assign MEM[12132] = MEM[338] + MEM[6465];
assign MEM[12133] = MEM[339] + MEM[5652];
assign MEM[12134] = MEM[340] + MEM[3237];
assign MEM[12135] = MEM[341] + MEM[5114];
assign MEM[12136] = MEM[343] + MEM[8380];
assign MEM[12137] = MEM[349] + MEM[10725];
assign MEM[12138] = MEM[354] + MEM[6206];
assign MEM[12139] = MEM[359] + MEM[6699];
assign MEM[12140] = MEM[363] + MEM[10660];
assign MEM[12141] = MEM[364] + MEM[6421];
assign MEM[12142] = MEM[365] + MEM[2670];
assign MEM[12143] = MEM[371] + MEM[2307];
assign MEM[12144] = MEM[373] + MEM[5052];
assign MEM[12145] = MEM[380] + MEM[1974];
assign MEM[12146] = MEM[381] + MEM[3924];
assign MEM[12147] = MEM[383] + MEM[3599];
assign MEM[12148] = MEM[387] + MEM[6054];
assign MEM[12149] = MEM[395] + MEM[4583];
assign MEM[12150] = MEM[398] + MEM[3058];
assign MEM[12151] = MEM[415] + MEM[7647];
assign MEM[12152] = MEM[422] + MEM[804];
assign MEM[12153] = MEM[429] + MEM[7448];
assign MEM[12154] = MEM[430] + MEM[3222];
assign MEM[12155] = MEM[431] + MEM[6629];
assign MEM[12156] = MEM[438] + MEM[3042];
assign MEM[12157] = MEM[445] + MEM[1427];
assign MEM[12158] = MEM[446] + MEM[4398];
assign MEM[12159] = MEM[447] + MEM[5167];
assign MEM[12160] = MEM[454] + MEM[9726];
assign MEM[12161] = MEM[455] + MEM[2406];
assign MEM[12162] = MEM[470] + MEM[6390];
assign MEM[12163] = MEM[471] + MEM[6888];
assign MEM[12164] = MEM[477] + MEM[8139];
assign MEM[12165] = MEM[483] + MEM[1111];
assign MEM[12166] = MEM[484] + MEM[7330];
assign MEM[12167] = MEM[487] + MEM[4783];
assign MEM[12168] = MEM[493] + MEM[1522];
assign MEM[12169] = MEM[495] + MEM[7730];
assign MEM[12170] = MEM[501] + MEM[10586];
assign MEM[12171] = MEM[507] + MEM[10605];
assign MEM[12172] = MEM[509] + MEM[4485];
assign MEM[12173] = MEM[514] + MEM[4886];
assign MEM[12174] = MEM[515] + MEM[1462];
assign MEM[12175] = MEM[517] + MEM[4522];
assign MEM[12176] = MEM[518] + MEM[31];
assign MEM[12177] = MEM[527] + MEM[5207];
assign MEM[12178] = MEM[530] + MEM[4251];
assign MEM[12179] = MEM[532] + MEM[4487];
assign MEM[12180] = MEM[534] + MEM[4391];
assign MEM[12181] = MEM[543] + MEM[5315];
assign MEM[12182] = MEM[547] + MEM[1863];
assign MEM[12183] = MEM[551] + MEM[3332];
assign MEM[12184] = MEM[554] + MEM[5035];
assign MEM[12185] = MEM[558] + MEM[2414];
assign MEM[12186] = MEM[559] + MEM[2046];
assign MEM[12187] = MEM[564] + MEM[8102];
assign MEM[12188] = MEM[566] + MEM[4866];
assign MEM[12189] = MEM[570] + MEM[693];
assign MEM[12190] = MEM[571] + MEM[7686];
assign MEM[12191] = MEM[574] + MEM[2324];
assign MEM[12192] = MEM[579] + MEM[2316];
assign MEM[12193] = MEM[586] + MEM[3891];
assign MEM[12194] = MEM[588] + MEM[4740];
assign MEM[12195] = MEM[591] + MEM[6111];
assign MEM[12196] = MEM[594] + MEM[6358];
assign MEM[12197] = MEM[596] + MEM[2051];
assign MEM[12198] = MEM[598] + MEM[5499];
assign MEM[12199] = MEM[602] + MEM[6123];
assign MEM[12200] = MEM[604] + MEM[1187];
assign MEM[12201] = MEM[607] + MEM[3837];
assign MEM[12202] = MEM[611] + MEM[727];
assign MEM[12203] = MEM[620] + MEM[6644];
assign MEM[12204] = MEM[621] + MEM[4228];
assign MEM[12205] = MEM[626] + MEM[2227];
assign MEM[12206] = MEM[627] + MEM[3108];
assign MEM[12207] = MEM[636] + MEM[6753];
assign MEM[12208] = MEM[639] + MEM[5915];
assign MEM[12209] = MEM[651] + MEM[1807];
assign MEM[12210] = MEM[652] + MEM[879];
assign MEM[12211] = MEM[653] + MEM[9315];
assign MEM[12212] = MEM[661] + MEM[1182];
assign MEM[12213] = MEM[663] + MEM[2508];
assign MEM[12214] = MEM[677] + MEM[10392];
assign MEM[12215] = MEM[678] + MEM[2181];
assign MEM[12216] = MEM[687] + MEM[8129];
assign MEM[12217] = MEM[695] + MEM[1716];
assign MEM[12218] = MEM[709] + MEM[1236];
assign MEM[12219] = MEM[711] + MEM[3189];
assign MEM[12220] = MEM[716] + MEM[2957];
assign MEM[12221] = MEM[723] + MEM[3030];
assign MEM[12222] = MEM[724] + MEM[3892];
assign MEM[12223] = MEM[730] + MEM[7106];
assign MEM[12224] = MEM[732] + MEM[2002];
assign MEM[12225] = MEM[733] + MEM[1436];
assign MEM[12226] = MEM[741] + MEM[7215];
assign MEM[12227] = MEM[758] + MEM[2595];
assign MEM[12228] = MEM[761] + MEM[1620];
assign MEM[12229] = MEM[765] + MEM[2788];
assign MEM[12230] = MEM[767] + MEM[3906];
assign MEM[12231] = MEM[771] + MEM[2023];
assign MEM[12232] = MEM[772] + MEM[1531];
assign MEM[12233] = MEM[774] + MEM[5787];
assign MEM[12234] = MEM[789] + MEM[764];
assign MEM[12235] = MEM[803] + MEM[5532];
assign MEM[12236] = MEM[812] + MEM[4023];
assign MEM[12237] = MEM[814] + MEM[3477];
assign MEM[12238] = MEM[820] + MEM[6698];
assign MEM[12239] = MEM[821] + MEM[3559];
assign MEM[12240] = MEM[827] + MEM[8085];
assign MEM[12241] = MEM[831] + MEM[1612];
assign MEM[12242] = MEM[834] + MEM[887];
assign MEM[12243] = MEM[836] + MEM[2015];
assign MEM[12244] = MEM[838] + MEM[4363];
assign MEM[12245] = MEM[850] + MEM[2437];
assign MEM[12246] = MEM[853] + MEM[910];
assign MEM[12247] = MEM[854] + MEM[7774];
assign MEM[12248] = MEM[859] + MEM[5046];
assign MEM[12249] = MEM[860] + MEM[4575];
assign MEM[12250] = MEM[861] + MEM[1874];
assign MEM[12251] = MEM[863] + MEM[3605];
assign MEM[12252] = MEM[878] + MEM[8178];
assign MEM[12253] = MEM[885] + MEM[525];
assign MEM[12254] = MEM[886] + MEM[5934];
assign MEM[12255] = MEM[893] + MEM[6878];
assign MEM[12256] = MEM[895] + MEM[4237];
assign MEM[12257] = MEM[911] + MEM[3877];
assign MEM[12258] = MEM[917] + MEM[3567];
assign MEM[12259] = MEM[925] + MEM[8038];
assign MEM[12260] = MEM[927] + MEM[10585];
assign MEM[12261] = MEM[932] + MEM[7294];
assign MEM[12262] = MEM[934] + MEM[5182];
assign MEM[12263] = MEM[940] + MEM[3613];
assign MEM[12264] = MEM[943] + MEM[9399];
assign MEM[12265] = MEM[946] + MEM[11005];
assign MEM[12266] = MEM[947] + MEM[1628];
assign MEM[12267] = MEM[949] + MEM[3604];
assign MEM[12268] = MEM[950] + MEM[4500];
assign MEM[12269] = MEM[957] + MEM[999];
assign MEM[12270] = MEM[958] + MEM[6306];
assign MEM[12271] = MEM[962] + MEM[7454];
assign MEM[12272] = MEM[964] + MEM[3646];
assign MEM[12273] = MEM[965] + MEM[2710];
assign MEM[12274] = MEM[974] + MEM[2140];
assign MEM[12275] = MEM[981] + MEM[655];
assign MEM[12276] = MEM[982] + MEM[3485];
assign MEM[12277] = MEM[983] + MEM[4644];
assign MEM[12278] = MEM[986] + MEM[4716];
assign MEM[12279] = MEM[987] + MEM[3514];
assign MEM[12280] = MEM[990] + MEM[407];
assign MEM[12281] = MEM[997] + MEM[4340];
assign MEM[12282] = MEM[1007] + MEM[7482];
assign MEM[12283] = MEM[1010] + MEM[3238];
assign MEM[12284] = MEM[1021] + MEM[4676];
assign MEM[12285] = MEM[1026] + MEM[2639];
assign MEM[12286] = MEM[1028] + MEM[1260];
assign MEM[12287] = MEM[1030] + MEM[2035];
assign MEM[12288] = MEM[1037] + MEM[2666];
assign MEM[12289] = MEM[1043] + MEM[1150];
assign MEM[12290] = MEM[1052] + MEM[2158];
assign MEM[12291] = MEM[1053] + MEM[1406];
assign MEM[12292] = MEM[1058] + MEM[2453];
assign MEM[12293] = MEM[1059] + MEM[1532];
assign MEM[12294] = MEM[1060] + MEM[2606];
assign MEM[12295] = MEM[1061] + MEM[1661];
assign MEM[12296] = MEM[1062] + MEM[2516];
assign MEM[12297] = MEM[1067] + MEM[5590];
assign MEM[12298] = MEM[1068] + MEM[1659];
assign MEM[12299] = MEM[1070] + MEM[1437];
assign MEM[12300] = MEM[1071] + MEM[5902];
assign MEM[12301] = MEM[1074] + MEM[9451];
assign MEM[12302] = MEM[1077] + MEM[1371];
assign MEM[12303] = MEM[1091] + MEM[2266];
assign MEM[12304] = MEM[1095] + MEM[6419];
assign MEM[12305] = MEM[1098] + MEM[5037];
assign MEM[12306] = MEM[1100] + MEM[3014];
assign MEM[12307] = MEM[1102] + MEM[1989];
assign MEM[12308] = MEM[1103] + MEM[1957];
assign MEM[12309] = MEM[1107] + MEM[406];
assign MEM[12310] = MEM[1109] + MEM[3707];
assign MEM[12311] = MEM[1110] + MEM[5981];
assign MEM[12312] = MEM[1117] + MEM[4498];
assign MEM[12313] = MEM[1119] + MEM[3554];
assign MEM[12314] = MEM[1126] + MEM[4738];
assign MEM[12315] = MEM[1135] + MEM[4239];
assign MEM[12316] = MEM[1142] + MEM[5092];
assign MEM[12317] = MEM[1148] + MEM[2879];
assign MEM[12318] = MEM[1151] + MEM[2399];
assign MEM[12319] = MEM[1155] + MEM[5451];
assign MEM[12320] = MEM[1156] + MEM[6156];
assign MEM[12321] = MEM[1158] + MEM[1739];
assign MEM[12322] = MEM[1159] + MEM[2950];
assign MEM[12323] = MEM[1163] + MEM[1443];
assign MEM[12324] = MEM[1164] + MEM[9376];
assign MEM[12325] = MEM[1165] + MEM[3660];
assign MEM[12326] = MEM[1166] + MEM[3843];
assign MEM[12327] = MEM[1171] + MEM[4645];
assign MEM[12328] = MEM[1175] + MEM[1748];
assign MEM[12329] = MEM[1178] + MEM[2038];
assign MEM[12330] = MEM[1180] + MEM[5642];
assign MEM[12331] = MEM[1190] + MEM[5421];
assign MEM[12332] = MEM[1195] + MEM[4347];
assign MEM[12333] = MEM[1197] + MEM[3156];
assign MEM[12334] = MEM[1198] + MEM[1574];
assign MEM[12335] = MEM[1202] + MEM[7261];
assign MEM[12336] = MEM[1211] + MEM[734];
assign MEM[12337] = MEM[1212] + MEM[1903];
assign MEM[12338] = MEM[1214] + MEM[2518];
assign MEM[12339] = MEM[1218] + MEM[1747];
assign MEM[12340] = MEM[1219] + MEM[4669];
assign MEM[12341] = MEM[1221] + MEM[1986];
assign MEM[12342] = MEM[1223] + MEM[3991];
assign MEM[12343] = MEM[1230] + MEM[2404];
assign MEM[12344] = MEM[1231] + MEM[10716];
assign MEM[12345] = MEM[1235] + MEM[1906];
assign MEM[12346] = MEM[1239] + MEM[10730];
assign MEM[12347] = MEM[1242] + MEM[4813];
assign MEM[12348] = MEM[1245] + MEM[3531];
assign MEM[12349] = MEM[1246] + MEM[5975];
assign MEM[12350] = MEM[1251] + MEM[8975];
assign MEM[12351] = MEM[1253] + MEM[5572];
assign MEM[12352] = MEM[1263] + MEM[1557];
assign MEM[12353] = MEM[1268] + MEM[2635];
assign MEM[12354] = MEM[1276] + MEM[2725];
assign MEM[12355] = MEM[1278] + MEM[6133];
assign MEM[12356] = MEM[1292] + MEM[2117];
assign MEM[12357] = MEM[1294] + MEM[2075];
assign MEM[12358] = MEM[1298] + MEM[3202];
assign MEM[12359] = MEM[1302] + MEM[531];
assign MEM[12360] = MEM[1308] + MEM[3471];
assign MEM[12361] = MEM[1309] + MEM[6895];
assign MEM[12362] = MEM[1315] + MEM[4556];
assign MEM[12363] = MEM[1322] + MEM[3213];
assign MEM[12364] = MEM[1324] + MEM[4511];
assign MEM[12365] = MEM[1327] + MEM[2563];
assign MEM[12366] = MEM[1332] + MEM[1587];
assign MEM[12367] = MEM[1333] + MEM[1565];
assign MEM[12368] = MEM[1334] + MEM[2187];
assign MEM[12369] = MEM[1335] + MEM[8511];
assign MEM[12370] = MEM[1342] + MEM[5643];
assign MEM[12371] = MEM[1349] + MEM[4972];
assign MEM[12372] = MEM[1374] + MEM[3375];
assign MEM[12373] = MEM[1375] + MEM[2740];
assign MEM[12374] = MEM[1380] + MEM[2014];
assign MEM[12375] = MEM[1381] + MEM[3166];
assign MEM[12376] = MEM[1387] + MEM[5428];
assign MEM[12377] = MEM[1389] + MEM[5645];
assign MEM[12378] = MEM[1390] + MEM[8061];
assign MEM[12379] = MEM[1396] + MEM[8391];
assign MEM[12380] = MEM[1397] + MEM[4754];
assign MEM[12381] = MEM[1398] + MEM[7581];
assign MEM[12382] = MEM[1404] + MEM[5012];
assign MEM[12383] = MEM[1405] + MEM[4387];
assign MEM[12384] = MEM[1407] + MEM[2558];
assign MEM[12385] = MEM[1410] + MEM[6729];
assign MEM[12386] = MEM[1411] + MEM[4692];
assign MEM[12387] = MEM[1414] + MEM[9322];
assign MEM[12388] = MEM[1420] + MEM[4906];
assign MEM[12389] = MEM[1422] + MEM[7790];
assign MEM[12390] = MEM[1423] + MEM[3879];
assign MEM[12391] = MEM[1429] + MEM[7483];
assign MEM[12392] = MEM[1438] + MEM[1900];
assign MEM[12393] = MEM[1439] + MEM[3611];
assign MEM[12394] = MEM[1444] + MEM[747];
assign MEM[12395] = MEM[1451] + MEM[4495];
assign MEM[12396] = MEM[1453] + MEM[1765];
assign MEM[12397] = MEM[1455] + MEM[5498];
assign MEM[12398] = MEM[1463] + MEM[4902];
assign MEM[12399] = MEM[1467] + MEM[4285];
assign MEM[12400] = MEM[1478] + MEM[2366];
assign MEM[12401] = MEM[1479] + MEM[1773];
assign MEM[12402] = MEM[1483] + MEM[6172];
assign MEM[12403] = MEM[1484] + MEM[6843];
assign MEM[12404] = MEM[1485] + MEM[3949];
assign MEM[12405] = MEM[1490] + MEM[1196];
assign MEM[12406] = MEM[1493] + MEM[3509];
assign MEM[12407] = MEM[1501] + MEM[6660];
assign MEM[12408] = MEM[1503] + MEM[6568];
assign MEM[12409] = MEM[1507] + MEM[3335];
assign MEM[12410] = MEM[1514] + MEM[2479];
assign MEM[12411] = MEM[1516] + MEM[7145];
assign MEM[12412] = MEM[1526] + MEM[2796];
assign MEM[12413] = MEM[1527] + MEM[5444];
assign MEM[12414] = MEM[1530] + MEM[3277];
assign MEM[12415] = MEM[1539] + MEM[4215];
assign MEM[12416] = MEM[1543] + MEM[5989];
assign MEM[12417] = MEM[1546] + MEM[4615];
assign MEM[12418] = MEM[1550] + MEM[2375];
assign MEM[12419] = MEM[1551] + MEM[5847];
assign MEM[12420] = MEM[1555] + MEM[2983];
assign MEM[12421] = MEM[1556] + MEM[622];
assign MEM[12422] = MEM[1563] + MEM[7721];
assign MEM[12423] = MEM[1564] + MEM[6324];
assign MEM[12424] = MEM[1566] + MEM[1734];
assign MEM[12425] = MEM[1578] + MEM[3884];
assign MEM[12426] = MEM[1579] + MEM[6155];
assign MEM[12427] = MEM[1583] + MEM[3630];
assign MEM[12428] = MEM[1594] + MEM[2127];
assign MEM[12429] = MEM[1595] + MEM[3290];
assign MEM[12430] = MEM[1598] + MEM[4075];
assign MEM[12431] = MEM[1599] + MEM[8513];
assign MEM[12432] = MEM[1603] + MEM[1862];
assign MEM[12433] = MEM[1604] + MEM[3383];
assign MEM[12434] = MEM[1605] + MEM[5942];
assign MEM[12435] = MEM[1615] + MEM[5462];
assign MEM[12436] = MEM[1618] + MEM[4950];
assign MEM[12437] = MEM[1619] + MEM[2564];
assign MEM[12438] = MEM[1626] + MEM[5186];
assign MEM[12439] = MEM[1629] + MEM[2931];
assign MEM[12440] = MEM[1630] + MEM[6473];
assign MEM[12441] = MEM[1636] + MEM[3162];
assign MEM[12442] = MEM[1637] + MEM[4082];
assign MEM[12443] = MEM[1638] + MEM[2372];
assign MEM[12444] = MEM[1646] + MEM[4283];
assign MEM[12445] = MEM[1647] + MEM[3461];
assign MEM[12446] = MEM[1650] + MEM[2847];
assign MEM[12447] = MEM[1652] + MEM[3708];
assign MEM[12448] = MEM[1653] + MEM[4415];
assign MEM[12449] = MEM[1655] + MEM[1134];
assign MEM[12450] = MEM[1668] + MEM[2383];
assign MEM[12451] = MEM[1671] + MEM[8495];
assign MEM[12452] = MEM[1678] + MEM[6857];
assign MEM[12453] = MEM[1679] + MEM[5962];
assign MEM[12454] = MEM[1685] + MEM[4164];
assign MEM[12455] = MEM[1686] + MEM[3639];
assign MEM[12456] = MEM[1687] + MEM[1700];
assign MEM[12457] = MEM[1692] + MEM[1972];
assign MEM[12458] = MEM[1702] + MEM[3948];
assign MEM[12459] = MEM[1707] + MEM[5519];
assign MEM[12460] = MEM[1715] + MEM[4159];
assign MEM[12461] = MEM[1723] + MEM[5948];
assign MEM[12462] = MEM[1727] + MEM[9028];
assign MEM[12463] = MEM[1732] + MEM[7828];
assign MEM[12464] = MEM[1735] + MEM[3652];
assign MEM[12465] = MEM[1740] + MEM[9099];
assign MEM[12466] = MEM[1742] + MEM[4155];
assign MEM[12467] = MEM[1743] + MEM[4797];
assign MEM[12468] = MEM[1751] + MEM[5322];
assign MEM[12469] = MEM[1758] + MEM[1982];
assign MEM[12470] = MEM[1764] + MEM[6047];
assign MEM[12471] = MEM[1767] + MEM[6675];
assign MEM[12472] = MEM[1771] + MEM[2478];
assign MEM[12473] = MEM[1779] + MEM[2028];
assign MEM[12474] = MEM[1783] + MEM[6614];
assign MEM[12475] = MEM[1789] + MEM[2484];
assign MEM[12476] = MEM[1791] + MEM[1838];
assign MEM[12477] = MEM[1803] + MEM[2709];
assign MEM[12478] = MEM[1804] + MEM[4639];
assign MEM[12479] = MEM[1814] + MEM[5463];
assign MEM[12480] = MEM[1815] + MEM[2491];
assign MEM[12481] = MEM[1822] + MEM[2498];
assign MEM[12482] = MEM[1829] + MEM[3740];
assign MEM[12483] = MEM[1839] + MEM[4579];
assign MEM[12484] = MEM[1843] + MEM[5575];
assign MEM[12485] = MEM[1845] + MEM[4686];
assign MEM[12486] = MEM[1851] + MEM[4292];
assign MEM[12487] = MEM[1853] + MEM[2767];
assign MEM[12488] = MEM[1854] + MEM[4524];
assign MEM[12489] = MEM[1859] + MEM[3405];
assign MEM[12490] = MEM[1868] + MEM[2468];
assign MEM[12491] = MEM[1870] + MEM[2863];
assign MEM[12492] = MEM[1875] + MEM[2511];
assign MEM[12493] = MEM[1876] + MEM[6061];
assign MEM[12494] = MEM[1877] + MEM[3538];
assign MEM[12495] = MEM[1878] + MEM[11038];
assign MEM[12496] = MEM[1887] + MEM[4318];
assign MEM[12497] = MEM[1893] + MEM[1970];
assign MEM[12498] = MEM[1894] + MEM[2135];
assign MEM[12499] = MEM[1899] + MEM[4430];
assign MEM[12500] = MEM[1901] + MEM[10903];
assign MEM[12501] = MEM[1907] + MEM[4820];
assign MEM[12502] = MEM[1908] + MEM[3823];
assign MEM[12503] = MEM[1909] + MEM[5699];
assign MEM[12504] = MEM[1910] + MEM[5717];
assign MEM[12505] = MEM[1911] + MEM[4324];
assign MEM[12506] = MEM[1916] + MEM[2502];
assign MEM[12507] = MEM[1918] + MEM[2142];
assign MEM[12508] = MEM[1919] + MEM[5628];
assign MEM[12509] = MEM[1923] + MEM[5534];
assign MEM[12510] = MEM[1926] + MEM[4762];
assign MEM[12511] = MEM[1934] + MEM[166];
assign MEM[12512] = MEM[1935] + MEM[2141];
assign MEM[12513] = MEM[1939] + MEM[10573];
assign MEM[12514] = MEM[1949] + MEM[4452];
assign MEM[12515] = MEM[1955] + MEM[6637];
assign MEM[12516] = MEM[1958] + MEM[3494];
assign MEM[12517] = MEM[1964] + MEM[5077];
assign MEM[12518] = MEM[1971] + MEM[5015];
assign MEM[12519] = MEM[1973] + MEM[8512];
assign MEM[12520] = MEM[1975] + MEM[1997];
assign MEM[12521] = MEM[1979] + MEM[7956];
assign MEM[12522] = MEM[1983] + MEM[2822];
assign MEM[12523] = MEM[1990] + MEM[6277];
assign MEM[12524] = MEM[1991] + MEM[10631];
assign MEM[12525] = MEM[1995] + MEM[4426];
assign MEM[12526] = MEM[2003] + MEM[7695];
assign MEM[12527] = MEM[2012] + MEM[2628];
assign MEM[12528] = MEM[2013] + MEM[7889];
assign MEM[12529] = MEM[2029] + MEM[3614];
assign MEM[12530] = MEM[2036] + MEM[7697];
assign MEM[12531] = MEM[2042] + MEM[3716];
assign MEM[12532] = MEM[2044] + MEM[4071];
assign MEM[12533] = MEM[2045] + MEM[8336];
assign MEM[12534] = MEM[2052] + MEM[6343];
assign MEM[12535] = MEM[2053] + MEM[10785];
assign MEM[12536] = MEM[2054] + MEM[6416];
assign MEM[12537] = MEM[2068] + MEM[3476];
assign MEM[12538] = MEM[2070] + MEM[5883];
assign MEM[12539] = MEM[2076] + MEM[3339];
assign MEM[12540] = MEM[2083] + MEM[703];
assign MEM[12541] = MEM[2085] + MEM[4566];
assign MEM[12542] = MEM[2093] + MEM[4261];
assign MEM[12543] = MEM[2095] + MEM[6389];
assign MEM[12544] = MEM[2098] + MEM[2268];
assign MEM[12545] = MEM[2107] + MEM[4658];
assign MEM[12546] = MEM[2110] + MEM[4910];
assign MEM[12547] = MEM[2115] + MEM[8477];
assign MEM[12548] = MEM[2116] + MEM[6007];
assign MEM[12549] = MEM[2122] + MEM[10208];
assign MEM[12550] = MEM[2124] + MEM[3314];
assign MEM[12551] = MEM[2126] + MEM[5111];
assign MEM[12552] = MEM[2132] + MEM[2221];
assign MEM[12553] = MEM[2147] + MEM[10609];
assign MEM[12554] = MEM[2148] + MEM[5399];
assign MEM[12555] = MEM[2155] + MEM[2830];
assign MEM[12556] = MEM[2157] + MEM[2974];
assign MEM[12557] = MEM[2163] + MEM[5351];
assign MEM[12558] = MEM[2167] + MEM[8095];
assign MEM[12559] = MEM[2172] + MEM[3895];
assign MEM[12560] = MEM[2174] + MEM[3667];
assign MEM[12561] = MEM[2179] + MEM[3683];
assign MEM[12562] = MEM[2183] + MEM[3157];
assign MEM[12563] = MEM[2190] + MEM[1607];
assign MEM[12564] = MEM[2196] + MEM[2538];
assign MEM[12565] = MEM[2204] + MEM[10667];
assign MEM[12566] = MEM[2211] + MEM[9292];
assign MEM[12567] = MEM[2214] + MEM[2267];
assign MEM[12568] = MEM[2219] + MEM[3828];
assign MEM[12569] = MEM[2223] + MEM[9334];
assign MEM[12570] = MEM[2228] + MEM[6887];
assign MEM[12571] = MEM[2229] + MEM[133];
assign MEM[12572] = MEM[2236] + MEM[1818];
assign MEM[12573] = MEM[2237] + MEM[10675];
assign MEM[12574] = MEM[2245] + MEM[7912];
assign MEM[12575] = MEM[2246] + MEM[3527];
assign MEM[12576] = MEM[2247] + MEM[4646];
assign MEM[12577] = MEM[2253] + MEM[5119];
assign MEM[12578] = MEM[2255] + MEM[6281];
assign MEM[12579] = MEM[2259] + MEM[3813];
assign MEM[12580] = MEM[2260] + MEM[6942];
assign MEM[12581] = MEM[2261] + MEM[3886];
assign MEM[12582] = MEM[2262] + MEM[5390];
assign MEM[12583] = MEM[2270] + MEM[3037];
assign MEM[12584] = MEM[2271] + MEM[8068];
assign MEM[12585] = MEM[2275] + MEM[7608];
assign MEM[12586] = MEM[2276] + MEM[2620];
assign MEM[12587] = MEM[2283] + MEM[4131];
assign MEM[12588] = MEM[2284] + MEM[2732];
assign MEM[12589] = MEM[2285] + MEM[7795];
assign MEM[12590] = MEM[2292] + MEM[877];
assign MEM[12591] = MEM[2303] + MEM[4540];
assign MEM[12592] = MEM[2306] + MEM[5469];
assign MEM[12593] = MEM[2310] + MEM[2566];
assign MEM[12594] = MEM[2314] + MEM[5359];
assign MEM[12595] = MEM[2318] + MEM[4973];
assign MEM[12596] = MEM[2319] + MEM[2701];
assign MEM[12597] = MEM[2322] + MEM[6367];
assign MEM[12598] = MEM[2330] + MEM[2373];
assign MEM[12599] = MEM[2332] + MEM[4867];
assign MEM[12600] = MEM[2341] + MEM[3379];
assign MEM[12601] = MEM[2342] + MEM[7114];
assign MEM[12602] = MEM[2343] + MEM[8533];
assign MEM[12603] = MEM[2350] + MEM[6715];
assign MEM[12604] = MEM[2357] + MEM[9889];
assign MEM[12605] = MEM[2358] + MEM[4436];
assign MEM[12606] = MEM[2362] + MEM[5669];
assign MEM[12607] = MEM[2363] + MEM[3628];
assign MEM[12608] = MEM[2370] + MEM[5260];
assign MEM[12609] = MEM[2371] + MEM[10726];
assign MEM[12610] = MEM[2380] + MEM[1445];
assign MEM[12611] = MEM[2381] + MEM[3204];
assign MEM[12612] = MEM[2382] + MEM[8544];
assign MEM[12613] = MEM[2390] + MEM[6853];
assign MEM[12614] = MEM[2391] + MEM[3111];
assign MEM[12615] = MEM[2394] + MEM[3436];
assign MEM[12616] = MEM[2396] + MEM[3474];
assign MEM[12617] = MEM[2398] + MEM[3005];
assign MEM[12618] = MEM[2402] + MEM[9383];
assign MEM[12619] = MEM[2405] + MEM[3731];
assign MEM[12620] = MEM[2407] + MEM[5685];
assign MEM[12621] = MEM[2411] + MEM[5589];
assign MEM[12622] = MEM[2412] + MEM[4406];
assign MEM[12623] = MEM[2418] + MEM[2531];
assign MEM[12624] = MEM[2420] + MEM[4439];
assign MEM[12625] = MEM[2429] + MEM[4778];
assign MEM[12626] = MEM[2430] + MEM[2991];
assign MEM[12627] = MEM[2435] + MEM[7902];
assign MEM[12628] = MEM[2439] + MEM[2891];
assign MEM[12629] = MEM[2443] + MEM[3051];
assign MEM[12630] = MEM[2445] + MEM[2845];
assign MEM[12631] = MEM[2446] + MEM[7974];
assign MEM[12632] = MEM[2450] + MEM[4743];
assign MEM[12633] = MEM[2460] + MEM[2846];
assign MEM[12634] = MEM[2469] + MEM[2903];
assign MEM[12635] = MEM[2471] + MEM[5211];
assign MEM[12636] = MEM[2476] + MEM[3475];
assign MEM[12637] = MEM[2493] + MEM[743];
assign MEM[12638] = MEM[2495] + MEM[173];
assign MEM[12639] = MEM[2506] + MEM[2758];
assign MEM[12640] = MEM[2509] + MEM[3763];
assign MEM[12641] = MEM[2532] + MEM[8080];
assign MEM[12642] = MEM[2533] + MEM[6297];
assign MEM[12643] = MEM[2540] + MEM[3226];
assign MEM[12644] = MEM[2543] + MEM[8656];
assign MEM[12645] = MEM[2548] + MEM[9054];
assign MEM[12646] = MEM[2549] + MEM[4621];
assign MEM[12647] = MEM[2565] + MEM[5788];
assign MEM[12648] = MEM[2572] + MEM[7849];
assign MEM[12649] = MEM[2573] + MEM[4890];
assign MEM[12650] = MEM[2575] + MEM[2813];
assign MEM[12651] = MEM[2580] + MEM[3979];
assign MEM[12652] = MEM[2587] + MEM[4091];
assign MEM[12653] = MEM[2591] + MEM[3291];
assign MEM[12654] = MEM[2594] + MEM[1186];
assign MEM[12655] = MEM[2596] + MEM[3212];
assign MEM[12656] = MEM[2597] + MEM[7744];
assign MEM[12657] = MEM[2615] + MEM[6069];
assign MEM[12658] = MEM[2621] + MEM[6739];
assign MEM[12659] = MEM[2626] + MEM[6329];
assign MEM[12660] = MEM[2627] + MEM[6746];
assign MEM[12661] = MEM[2634] + MEM[8122];
assign MEM[12662] = MEM[2636] + MEM[4631];
assign MEM[12663] = MEM[2638] + MEM[7430];
assign MEM[12664] = MEM[2643] + MEM[3699];
assign MEM[12665] = MEM[2650] + MEM[5738];
assign MEM[12666] = MEM[2654] + MEM[3295];
assign MEM[12667] = MEM[2663] + MEM[10776];
assign MEM[12668] = MEM[2676] + MEM[4319];
assign MEM[12669] = MEM[2687] + MEM[742];
assign MEM[12670] = MEM[2702] + MEM[5347];
assign MEM[12671] = MEM[2706] + MEM[5013];
assign MEM[12672] = MEM[2714] + MEM[7440];
assign MEM[12673] = MEM[2719] + MEM[1509];
assign MEM[12674] = MEM[2724] + MEM[6745];
assign MEM[12675] = MEM[2731] + MEM[3523];
assign MEM[12676] = MEM[2735] + MEM[7726];
assign MEM[12677] = MEM[2742] + MEM[3930];
assign MEM[12678] = MEM[2751] + MEM[3966];
assign MEM[12679] = MEM[2755] + MEM[4806];
assign MEM[12680] = MEM[2756] + MEM[3331];
assign MEM[12681] = MEM[2764] + MEM[3706];
assign MEM[12682] = MEM[2770] + MEM[3271];
assign MEM[12683] = MEM[2778] + MEM[8076];
assign MEM[12684] = MEM[2779] + MEM[4654];
assign MEM[12685] = MEM[2782] + MEM[4165];
assign MEM[12686] = MEM[2790] + MEM[3230];
assign MEM[12687] = MEM[2794] + MEM[9081];
assign MEM[12688] = MEM[2798] + MEM[1039];
assign MEM[12689] = MEM[2799] + MEM[4029];
assign MEM[12690] = MEM[2807] + MEM[6287];
assign MEM[12691] = MEM[2815] + MEM[10466];
assign MEM[12692] = MEM[2820] + MEM[5551];
assign MEM[12693] = MEM[2842] + MEM[4431];
assign MEM[12694] = MEM[2851] + MEM[6812];
assign MEM[12695] = MEM[2858] + MEM[5533];
assign MEM[12696] = MEM[2861] + MEM[2919];
assign MEM[12697] = MEM[2862] + MEM[5691];
assign MEM[12698] = MEM[2869] + MEM[8504];
assign MEM[12699] = MEM[2886] + MEM[7091];
assign MEM[12700] = MEM[2887] + MEM[6584];
assign MEM[12701] = MEM[2892] + MEM[3756];
assign MEM[12702] = MEM[2909] + MEM[4238];
assign MEM[12703] = MEM[2911] + MEM[5477];
assign MEM[12704] = MEM[2926] + MEM[6775];
assign MEM[12705] = MEM[2933] + MEM[5431];
assign MEM[12706] = MEM[2934] + MEM[7256];
assign MEM[12707] = MEM[2935] + MEM[3445];
assign MEM[12708] = MEM[2949] + MEM[9631];
assign MEM[12709] = MEM[2955] + MEM[3063];
assign MEM[12710] = MEM[2956] + MEM[7328];
assign MEM[12711] = MEM[2967] + MEM[3590];
assign MEM[12712] = MEM[2995] + MEM[9067];
assign MEM[12713] = MEM[2999] + MEM[3915];
assign MEM[12714] = MEM[3004] + MEM[7983];
assign MEM[12715] = MEM[3006] + MEM[9367];
assign MEM[12716] = MEM[3010] + MEM[7668];
assign MEM[12717] = MEM[3015] + MEM[3197];
assign MEM[12718] = MEM[3022] + MEM[2378];
assign MEM[12719] = MEM[3039] + MEM[8927];
assign MEM[12720] = MEM[3043] + MEM[3490];
assign MEM[12721] = MEM[3045] + MEM[3207];
assign MEM[12722] = MEM[3055] + MEM[3622];
assign MEM[12723] = MEM[3059] + MEM[1684];
assign MEM[12724] = MEM[3068] + MEM[4770];
assign MEM[12725] = MEM[3069] + MEM[3453];
assign MEM[12726] = MEM[3075] + MEM[3943];
assign MEM[12727] = MEM[3094] + MEM[3359];
assign MEM[12728] = MEM[3100] + MEM[4287];
assign MEM[12729] = MEM[3103] + MEM[3292];
assign MEM[12730] = MEM[3114] + MEM[7511];
assign MEM[12731] = MEM[3115] + MEM[5892];
assign MEM[12732] = MEM[3118] + MEM[2941];
assign MEM[12733] = MEM[3119] + MEM[5415];
assign MEM[12734] = MEM[3127] + MEM[4246];
assign MEM[12735] = MEM[3132] + MEM[4206];
assign MEM[12736] = MEM[3151] + MEM[3287];
assign MEM[12737] = MEM[3170] + MEM[3733];
assign MEM[12738] = MEM[3174] + MEM[10445];
assign MEM[12739] = MEM[3185] + MEM[8489];
assign MEM[12740] = MEM[3190] + MEM[4747];
assign MEM[12741] = MEM[3191] + MEM[5634];
assign MEM[12742] = MEM[3195] + MEM[1895];
assign MEM[12743] = MEM[3196] + MEM[8260];
assign MEM[12744] = MEM[3198] + MEM[2677];
assign MEM[12745] = MEM[3205] + MEM[4059];
assign MEM[12746] = MEM[3206] + MEM[7489];
assign MEM[12747] = MEM[3210] + MEM[4213];
assign MEM[12748] = MEM[3211] + MEM[3621];
assign MEM[12749] = MEM[3227] + MEM[6486];
assign MEM[12750] = MEM[3231] + MEM[10697];
assign MEM[12751] = MEM[3236] + MEM[4829];
assign MEM[12752] = MEM[3243] + MEM[4967];
assign MEM[12753] = MEM[3246] + MEM[7003];
assign MEM[12754] = MEM[3251] + MEM[8583];
assign MEM[12755] = MEM[3252] + MEM[7568];
assign MEM[12756] = MEM[3259] + MEM[4494];
assign MEM[12757] = MEM[3260] + MEM[6755];
assign MEM[12758] = MEM[3262] + MEM[6983];
assign MEM[12759] = MEM[3269] + MEM[3502];
assign MEM[12760] = MEM[3275] + MEM[2111];
assign MEM[12761] = MEM[3283] + MEM[4735];
assign MEM[12762] = MEM[3294] + MEM[4348];
assign MEM[12763] = MEM[3308] + MEM[5285];
assign MEM[12764] = MEM[3317] + MEM[7818];
assign MEM[12765] = MEM[3318] + MEM[5567];
assign MEM[12766] = MEM[3319] + MEM[4997];
assign MEM[12767] = MEM[3324] + MEM[9045];
assign MEM[12768] = MEM[3330] + MEM[4196];
assign MEM[12769] = MEM[3333] + MEM[8263];
assign MEM[12770] = MEM[3338] + MEM[7211];
assign MEM[12771] = MEM[3348] + MEM[7011];
assign MEM[12772] = MEM[3350] + MEM[5591];
assign MEM[12773] = MEM[3371] + MEM[4157];
assign MEM[12774] = MEM[3374] + MEM[4683];
assign MEM[12775] = MEM[3380] + MEM[963];
assign MEM[12776] = MEM[3381] + MEM[4638];
assign MEM[12777] = MEM[3387] + MEM[8643];
assign MEM[12778] = MEM[3391] + MEM[7519];
assign MEM[12779] = MEM[3394] + MEM[7180];
assign MEM[12780] = MEM[3398] + MEM[4375];
assign MEM[12781] = MEM[3411] + MEM[7749];
assign MEM[12782] = MEM[3419] + MEM[4322];
assign MEM[12783] = MEM[3421] + MEM[6907];
assign MEM[12784] = MEM[3430] + MEM[10582];
assign MEM[12785] = MEM[3434] + MEM[3487];
assign MEM[12786] = MEM[3444] + MEM[6517];
assign MEM[12787] = MEM[3452] + MEM[4399];
assign MEM[12788] = MEM[3454] + MEM[1460];
assign MEM[12789] = MEM[3458] + MEM[4812];
assign MEM[12790] = MEM[3462] + MEM[6558];
assign MEM[12791] = MEM[3467] + MEM[8792];
assign MEM[12792] = MEM[3478] + MEM[3999];
assign MEM[12793] = MEM[3484] + MEM[7083];
assign MEM[12794] = MEM[3499] + MEM[3678];
assign MEM[12795] = MEM[3503] + MEM[2131];
assign MEM[12796] = MEM[3507] + MEM[5262];
assign MEM[12797] = MEM[3508] + MEM[4333];
assign MEM[12798] = MEM[3511] + MEM[7104];
assign MEM[12799] = MEM[3515] + MEM[3982];
assign MEM[12800] = MEM[3516] + MEM[3546];
assign MEM[12801] = MEM[3525] + MEM[7177];
assign MEM[12802] = MEM[3539] + MEM[3973];
assign MEM[12803] = MEM[3547] + MEM[2943];
assign MEM[12804] = MEM[3558] + MEM[7107];
assign MEM[12805] = MEM[3562] + MEM[1998];
assign MEM[12806] = MEM[3563] + MEM[5491];
assign MEM[12807] = MEM[3570] + MEM[4508];
assign MEM[12808] = MEM[3572] + MEM[10476];
assign MEM[12809] = MEM[3575] + MEM[4343];
assign MEM[12810] = MEM[3581] + MEM[6189];
assign MEM[12811] = MEM[3583] + MEM[9158];
assign MEM[12812] = MEM[3591] + MEM[1710];
assign MEM[12813] = MEM[3602] + MEM[8961];
assign MEM[12814] = MEM[3607] + MEM[7932];
assign MEM[12815] = MEM[3627] + MEM[7617];
assign MEM[12816] = MEM[3635] + MEM[3650];
assign MEM[12817] = MEM[3637] + MEM[10590];
assign MEM[12818] = MEM[3638] + MEM[3858];
assign MEM[12819] = MEM[3663] + MEM[4799];
assign MEM[12820] = MEM[3669] + MEM[9900];
assign MEM[12821] = MEM[3670] + MEM[3935];
assign MEM[12822] = MEM[3686] + MEM[6754];
assign MEM[12823] = MEM[3690] + MEM[3778];
assign MEM[12824] = MEM[3694] + MEM[10861];
assign MEM[12825] = MEM[3695] + MEM[5183];
assign MEM[12826] = MEM[3702] + MEM[5291];
assign MEM[12827] = MEM[3709] + MEM[5446];
assign MEM[12828] = MEM[3726] + MEM[5484];
assign MEM[12829] = MEM[3727] + MEM[6847];
assign MEM[12830] = MEM[3741] + MEM[4115];
assign MEM[12831] = MEM[3742] + MEM[2239];
assign MEM[12832] = MEM[3746] + MEM[6608];
assign MEM[12833] = MEM[3748] + MEM[7155];
assign MEM[12834] = MEM[3749] + MEM[4790];
assign MEM[12835] = MEM[3755] + MEM[762];
assign MEM[12836] = MEM[3762] + MEM[11092];
assign MEM[12837] = MEM[3766] + MEM[8147];
assign MEM[12838] = MEM[3770] + MEM[7559];
assign MEM[12839] = MEM[3772] + MEM[8744];
assign MEM[12840] = MEM[3774] + MEM[5301];
assign MEM[12841] = MEM[3779] + MEM[4623];
assign MEM[12842] = MEM[3789] + MEM[7465];
assign MEM[12843] = MEM[3795] + MEM[4204];
assign MEM[12844] = MEM[3798] + MEM[954];
assign MEM[12845] = MEM[3799] + MEM[6455];
assign MEM[12846] = MEM[3804] + MEM[5887];
assign MEM[12847] = MEM[3822] + MEM[10598];
assign MEM[12848] = MEM[3831] + MEM[3875];
assign MEM[12849] = MEM[3836] + MEM[7980];
assign MEM[12850] = MEM[3838] + MEM[4670];
assign MEM[12851] = MEM[3846] + MEM[6877];
assign MEM[12852] = MEM[3853] + MEM[4460];
assign MEM[12853] = MEM[3854] + MEM[7137];
assign MEM[12854] = MEM[3862] + MEM[5878];
assign MEM[12855] = MEM[3863] + MEM[4156];
assign MEM[12856] = MEM[3885] + MEM[6269];
assign MEM[12857] = MEM[3893] + MEM[8993];
assign MEM[12858] = MEM[3898] + MEM[7884];
assign MEM[12859] = MEM[3911] + MEM[6846];
assign MEM[12860] = MEM[3923] + MEM[6984];
assign MEM[12861] = MEM[3933] + MEM[4326];
assign MEM[12862] = MEM[3940] + MEM[2684];
assign MEM[12863] = MEM[3942] + MEM[10635];
assign MEM[12864] = MEM[3946] + MEM[5340];
assign MEM[12865] = MEM[3956] + MEM[8121];
assign MEM[12866] = MEM[3958] + MEM[4051];
assign MEM[12867] = MEM[3964] + MEM[4086];
assign MEM[12868] = MEM[3965] + MEM[7692];
assign MEM[12869] = MEM[3978] + MEM[2134];
assign MEM[12870] = MEM[3988] + MEM[7291];
assign MEM[12871] = MEM[3989] + MEM[5722];
assign MEM[12872] = MEM[3996] + MEM[4733];
assign MEM[12873] = MEM[4002] + MEM[5731];
assign MEM[12874] = MEM[4006] + MEM[6569];
assign MEM[12875] = MEM[4011] + MEM[4787];
assign MEM[12876] = MEM[4012] + MEM[6580];
assign MEM[12877] = MEM[4015] + MEM[5899];
assign MEM[12878] = MEM[4018] + MEM[9071];
assign MEM[12879] = MEM[4022] + MEM[8953];
assign MEM[12880] = MEM[4037] + MEM[6335];
assign MEM[12881] = MEM[4052] + MEM[6682];
assign MEM[12882] = MEM[4053] + MEM[9510];
assign MEM[12883] = MEM[4060] + MEM[6376];
assign MEM[12884] = MEM[4062] + MEM[10612];
assign MEM[12885] = MEM[4067] + MEM[6003];
assign MEM[12886] = MEM[4069] + MEM[7920];
assign MEM[12887] = MEM[4076] + MEM[4501];
assign MEM[12888] = MEM[4078] + MEM[1508];
assign MEM[12889] = MEM[4079] + MEM[5558];
assign MEM[12890] = MEM[4083] + MEM[7866];
assign MEM[12891] = MEM[4087] + MEM[5783];
assign MEM[12892] = MEM[4092] + MEM[7351];
assign MEM[12893] = MEM[4093] + MEM[966];
assign MEM[12894] = MEM[4095] + MEM[7917];
assign MEM[12895] = MEM[4098] + MEM[8075];
assign MEM[12896] = MEM[4099] + MEM[6174];
assign MEM[12897] = MEM[4102] + MEM[7966];
assign MEM[12898] = MEM[4106] + MEM[10639];
assign MEM[12899] = MEM[4108] + MEM[2364];
assign MEM[12900] = MEM[4110] + MEM[4132];
assign MEM[12901] = MEM[4111] + MEM[2653];
assign MEM[12902] = MEM[4114] + MEM[8096];
assign MEM[12903] = MEM[4116] + MEM[5736];
assign MEM[12904] = MEM[4118] + MEM[10856];
assign MEM[12905] = MEM[4122] + MEM[7516];
assign MEM[12906] = MEM[4126] + MEM[5229];
assign MEM[12907] = MEM[4139] + MEM[7708];
assign MEM[12908] = MEM[4140] + MEM[7332];
assign MEM[12909] = MEM[4143] + MEM[5006];
assign MEM[12910] = MEM[4149] + MEM[6670];
assign MEM[12911] = MEM[4158] + MEM[4191];
assign MEM[12912] = MEM[4166] + MEM[8713];
assign MEM[12913] = MEM[4173] + MEM[5252];
assign MEM[12914] = MEM[4174] + MEM[9052];
assign MEM[12915] = MEM[4186] + MEM[7122];
assign MEM[12916] = MEM[4188] + MEM[1749];
assign MEM[12917] = MEM[4189] + MEM[9422];
assign MEM[12918] = MEM[4205] + MEM[9171];
assign MEM[12919] = MEM[4207] + MEM[9240];
assign MEM[12920] = MEM[4211] + MEM[6903];
assign MEM[12921] = MEM[4218] + MEM[9153];
assign MEM[12922] = MEM[4220] + MEM[9130];
assign MEM[12923] = MEM[4221] + MEM[8015];
assign MEM[12924] = MEM[4223] + MEM[4884];
assign MEM[12925] = MEM[4231] + MEM[5538];
assign MEM[12926] = MEM[4245] + MEM[5243];
assign MEM[12927] = MEM[4247] + MEM[7285];
assign MEM[12928] = MEM[4255] + MEM[7340];
assign MEM[12929] = MEM[4271] + MEM[6154];
assign MEM[12930] = MEM[4282] + MEM[3972];
assign MEM[12931] = MEM[4291] + MEM[7592];
assign MEM[12932] = MEM[4293] + MEM[6923];
assign MEM[12933] = MEM[4295] + MEM[4335];
assign MEM[12934] = MEM[4298] + MEM[10808];
assign MEM[12935] = MEM[4303] + MEM[6166];
assign MEM[12936] = MEM[4307] + MEM[8081];
assign MEM[12937] = MEM[4308] + MEM[5905];
assign MEM[12938] = MEM[4314] + MEM[4926];
assign MEM[12939] = MEM[4317] + MEM[6678];
assign MEM[12940] = MEM[4327] + MEM[10591];
assign MEM[12941] = MEM[4338] + MEM[6262];
assign MEM[12942] = MEM[4341] + MEM[5143];
assign MEM[12943] = MEM[4346] + MEM[7610];
assign MEM[12944] = MEM[4349] + MEM[8979];
assign MEM[12945] = MEM[4355] + MEM[5741];
assign MEM[12946] = MEM[4357] + MEM[5341];
assign MEM[12947] = MEM[4365] + MEM[5631];
assign MEM[12948] = MEM[4367] + MEM[8091];
assign MEM[12949] = MEM[4383] + MEM[10545];
assign MEM[12950] = MEM[4407] + MEM[4717];
assign MEM[12951] = MEM[4412] + MEM[6142];
assign MEM[12952] = MEM[4413] + MEM[1810];
assign MEM[12953] = MEM[4420] + MEM[6116];
assign MEM[12954] = MEM[4423] + MEM[6290];
assign MEM[12955] = MEM[4435] + MEM[5076];
assign MEM[12956] = MEM[4437] + MEM[5829];
assign MEM[12957] = MEM[4443] + MEM[4839];
assign MEM[12958] = MEM[4446] + MEM[4674];
assign MEM[12959] = MEM[4451] + MEM[7615];
assign MEM[12960] = MEM[4466] + MEM[7810];
assign MEM[12961] = MEM[4469] + MEM[7203];
assign MEM[12962] = MEM[4470] + MEM[7311];
assign MEM[12963] = MEM[4477] + MEM[10951];
assign MEM[12964] = MEM[4478] + MEM[4558];
assign MEM[12965] = MEM[4493] + MEM[7672];
assign MEM[12966] = MEM[4502] + MEM[3730];
assign MEM[12967] = MEM[4506] + MEM[6560];
assign MEM[12968] = MEM[4509] + MEM[5492];
assign MEM[12969] = MEM[4530] + MEM[9879];
assign MEM[12970] = MEM[4532] + MEM[6537];
assign MEM[12971] = MEM[4546] + MEM[5703];
assign MEM[12972] = MEM[4548] + MEM[5813];
assign MEM[12973] = MEM[4550] + MEM[5918];
assign MEM[12974] = MEM[4559] + MEM[5766];
assign MEM[12975] = MEM[4563] + MEM[3806];
assign MEM[12976] = MEM[4564] + MEM[5959];
assign MEM[12977] = MEM[4567] + MEM[7977];
assign MEM[12978] = MEM[4571] + MEM[10834];
assign MEM[12979] = MEM[4572] + MEM[5506];
assign MEM[12980] = MEM[4574] + MEM[1675];
assign MEM[12981] = MEM[4581] + MEM[10705];
assign MEM[12982] = MEM[4582] + MEM[5227];
assign MEM[12983] = MEM[4587] + MEM[5781];
assign MEM[12984] = MEM[4591] + MEM[10678];
assign MEM[12985] = MEM[4597] + MEM[8902];
assign MEM[12986] = MEM[4598] + MEM[6940];
assign MEM[12987] = MEM[4604] + MEM[7154];
assign MEM[12988] = MEM[4611] + MEM[10820];
assign MEM[12989] = MEM[4612] + MEM[4883];
assign MEM[12990] = MEM[4613] + MEM[8175];
assign MEM[12991] = MEM[4614] + MEM[5636];
assign MEM[12992] = MEM[4619] + MEM[9757];
assign MEM[12993] = MEM[4620] + MEM[4450];
assign MEM[12994] = MEM[4647] + MEM[3659];
assign MEM[12995] = MEM[4650] + MEM[5646];
assign MEM[12996] = MEM[4653] + MEM[6706];
assign MEM[12997] = MEM[4666] + MEM[6725];
assign MEM[12998] = MEM[4671] + MEM[10616];
assign MEM[12999] = MEM[4675] + MEM[1927];
assign MEM[13000] = MEM[4685] + MEM[5890];
assign MEM[13001] = MEM[4709] + MEM[7123];
assign MEM[13002] = MEM[4711] + MEM[5879];
assign MEM[13003] = MEM[4715] + MEM[5906];
assign MEM[13004] = MEM[4722] + MEM[5397];
assign MEM[13005] = MEM[4723] + MEM[8590];
assign MEM[13006] = MEM[4724] + MEM[4781];
assign MEM[13007] = MEM[4725] + MEM[4148];
assign MEM[13008] = MEM[4727] + MEM[7613];
assign MEM[13009] = MEM[4730] + MEM[5330];
assign MEM[13010] = MEM[4748] + MEM[1943];
assign MEM[13011] = MEM[4751] + MEM[5494];
assign MEM[13012] = MEM[4766] + MEM[5036];
assign MEM[13013] = MEM[4782] + MEM[5667];
assign MEM[13014] = MEM[4788] + MEM[6849];
assign MEM[13015] = MEM[4794] + MEM[5418];
assign MEM[13016] = MEM[4796] + MEM[5435];
assign MEM[13017] = MEM[4798] + MEM[3323];
assign MEM[13018] = MEM[4811] + MEM[4942];
assign MEM[13019] = MEM[4818] + MEM[6901];
assign MEM[13020] = MEM[4821] + MEM[7365];
assign MEM[13021] = MEM[4822] + MEM[8376];
assign MEM[13022] = MEM[4828] + MEM[6430];
assign MEM[13023] = MEM[4830] + MEM[5075];
assign MEM[13024] = MEM[4836] + MEM[10175];
assign MEM[13025] = MEM[4843] + MEM[1469];
assign MEM[13026] = MEM[4844] + MEM[6921];
assign MEM[13027] = MEM[4845] + MEM[7967];
assign MEM[13028] = MEM[4862] + MEM[10997];
assign MEM[13029] = MEM[4870] + MEM[4605];
assign MEM[13030] = MEM[4871] + MEM[7481];
assign MEM[13031] = MEM[4874] + MEM[538];
assign MEM[13032] = MEM[4875] + MEM[7537];
assign MEM[13033] = MEM[4876] + MEM[2138];
assign MEM[13034] = MEM[4877] + MEM[5566];
assign MEM[13035] = MEM[4879] + MEM[9029];
assign MEM[13036] = MEM[4895] + MEM[5085];
assign MEM[13037] = MEM[4900] + MEM[9089];
assign MEM[13038] = MEM[4901] + MEM[6270];
assign MEM[13039] = MEM[4903] + MEM[8691];
assign MEM[13040] = MEM[4908] + MEM[5381];
assign MEM[13041] = MEM[4916] + MEM[6440];
assign MEM[13042] = MEM[4917] + MEM[7614];
assign MEM[13043] = MEM[4918] + MEM[6570];
assign MEM[13044] = MEM[4919] + MEM[6203];
assign MEM[13045] = MEM[4933] + MEM[7838];
assign MEM[13046] = MEM[4947] + MEM[5239];
assign MEM[13047] = MEM[4948] + MEM[5021];
assign MEM[13048] = MEM[4954] + MEM[7153];
assign MEM[13049] = MEM[4959] + MEM[7623];
assign MEM[13050] = MEM[4966] + MEM[5746];
assign MEM[13051] = MEM[4975] + MEM[5235];
assign MEM[13052] = MEM[4981] + MEM[5468];
assign MEM[13053] = MEM[4983] + MEM[7803];
assign MEM[13054] = MEM[4988] + MEM[7574];
assign MEM[13055] = MEM[4999] + MEM[7688];
assign MEM[13056] = MEM[5004] + MEM[10606];
assign MEM[13057] = MEM[5007] + MEM[3131];
assign MEM[13058] = MEM[5028] + MEM[5234];
assign MEM[13059] = MEM[5029] + MEM[3310];
assign MEM[13060] = MEM[5039] + MEM[5287];
assign MEM[13061] = MEM[5044] + MEM[5045];
assign MEM[13062] = MEM[5047] + MEM[6046];
assign MEM[13063] = MEM[5053] + MEM[6426];
assign MEM[13064] = MEM[5059] + MEM[5179];
assign MEM[13065] = MEM[5062] + MEM[6586];
assign MEM[13066] = MEM[5063] + MEM[6514];
assign MEM[13067] = MEM[5071] + MEM[8252];
assign MEM[13068] = MEM[5079] + MEM[10638];
assign MEM[13069] = MEM[5093] + MEM[5922];
assign MEM[13070] = MEM[5094] + MEM[9443];
assign MEM[13071] = MEM[5099] + MEM[6435];
assign MEM[13072] = MEM[5102] + MEM[1756];
assign MEM[13073] = MEM[5115] + MEM[4127];
assign MEM[13074] = MEM[5116] + MEM[8485];
assign MEM[13075] = MEM[5117] + MEM[5413];
assign MEM[13076] = MEM[5123] + MEM[5861];
assign MEM[13077] = MEM[5127] + MEM[6738];
assign MEM[13078] = MEM[5134] + MEM[5335];
assign MEM[13079] = MEM[5141] + MEM[5644];
assign MEM[13080] = MEM[5159] + MEM[10773];
assign MEM[13081] = MEM[5178] + MEM[5579];
assign MEM[13082] = MEM[5187] + MEM[7599];
assign MEM[13083] = MEM[5188] + MEM[7579];
assign MEM[13084] = MEM[5191] + MEM[6619];
assign MEM[13085] = MEM[5194] + MEM[7373];
assign MEM[13086] = MEM[5196] + MEM[1596];
assign MEM[13087] = MEM[5199] + MEM[7580];
assign MEM[13088] = MEM[5203] + MEM[1066];
assign MEM[13089] = MEM[5213] + MEM[7713];
assign MEM[13090] = MEM[5214] + MEM[3548];
assign MEM[13091] = MEM[5220] + MEM[9478];
assign MEM[13092] = MEM[5223] + MEM[8113];
assign MEM[13093] = MEM[5228] + MEM[978];
assign MEM[13094] = MEM[5244] + MEM[7957];
assign MEM[13095] = MEM[5245] + MEM[7797];
assign MEM[13096] = MEM[5253] + MEM[7995];
assign MEM[13097] = MEM[5261] + MEM[7225];
assign MEM[13098] = MEM[5263] + MEM[11295];
assign MEM[13099] = MEM[5266] + MEM[8101];
assign MEM[13100] = MEM[5269] + MEM[10771];
assign MEM[13101] = MEM[5270] + MEM[6536];
assign MEM[13102] = MEM[5278] + MEM[4907];
assign MEM[13103] = MEM[5279] + MEM[10810];
assign MEM[13104] = MEM[5283] + MEM[7414];
assign MEM[13105] = MEM[5284] + MEM[2286];
assign MEM[13106] = MEM[5292] + MEM[1891];
assign MEM[13107] = MEM[5294] + MEM[10151];
assign MEM[13108] = MEM[5295] + MEM[9114];
assign MEM[13109] = MEM[5299] + MEM[6703];
assign MEM[13110] = MEM[5302] + MEM[3860];
assign MEM[13111] = MEM[5303] + MEM[6532];
assign MEM[13112] = MEM[5314] + MEM[9468];
assign MEM[13113] = MEM[5316] + MEM[6354];
assign MEM[13114] = MEM[5318] + MEM[8911];
assign MEM[13115] = MEM[5319] + MEM[7350];
assign MEM[13116] = MEM[5325] + MEM[6917];
assign MEM[13117] = MEM[5331] + MEM[8571];
assign MEM[13118] = MEM[5334] + MEM[10812];
assign MEM[13119] = MEM[5343] + MEM[1500];
assign MEM[13120] = MEM[5366] + MEM[4499];
assign MEM[13121] = MEM[5367] + MEM[10685];
assign MEM[13122] = MEM[5382] + MEM[5718];
assign MEM[13123] = MEM[5391] + MEM[1063];
assign MEM[13124] = MEM[5404] + MEM[6611];
assign MEM[13125] = MEM[5405] + MEM[5445];
assign MEM[13126] = MEM[5406] + MEM[10749];
assign MEM[13127] = MEM[5411] + MEM[7282];
assign MEM[13128] = MEM[5419] + MEM[5524];
assign MEM[13129] = MEM[5423] + MEM[10768];
assign MEM[13130] = MEM[5439] + MEM[3629];
assign MEM[13131] = MEM[5442] + MEM[2853];
assign MEM[13132] = MEM[5447] + MEM[8290];
assign MEM[13133] = MEM[5452] + MEM[3279];
assign MEM[13134] = MEM[5453] + MEM[2550];
assign MEM[13135] = MEM[5454] + MEM[5502];
assign MEM[13136] = MEM[5458] + MEM[6801];
assign MEM[13137] = MEM[5475] + MEM[8236];
assign MEM[13138] = MEM[5476] + MEM[7043];
assign MEM[13139] = MEM[5483] + MEM[5997];
assign MEM[13140] = MEM[5500] + MEM[2996];
assign MEM[13141] = MEM[5501] + MEM[331];
assign MEM[13142] = MEM[5509] + MEM[8400];
assign MEM[13143] = MEM[5511] + MEM[2317];
assign MEM[13144] = MEM[5516] + MEM[5084];
assign MEM[13145] = MEM[5517] + MEM[6474];
assign MEM[13146] = MEM[5522] + MEM[8608];
assign MEM[13147] = MEM[5523] + MEM[6162];
assign MEM[13148] = MEM[5526] + MEM[5937];
assign MEM[13149] = MEM[5530] + MEM[8916];
assign MEM[13150] = MEM[5546] + MEM[3486];
assign MEM[13151] = MEM[5547] + MEM[7691];
assign MEM[13152] = MEM[5554] + MEM[8149];
assign MEM[13153] = MEM[5555] + MEM[10580];
assign MEM[13154] = MEM[5556] + MEM[3483];
assign MEM[13155] = MEM[5563] + MEM[4763];
assign MEM[13156] = MEM[5564] + MEM[10581];
assign MEM[13157] = MEM[5565] + MEM[2199];
assign MEM[13158] = MEM[5570] + MEM[10718];
assign MEM[13159] = MEM[5574] + MEM[3219];
assign MEM[13160] = MEM[5581] + MEM[5663];
assign MEM[13161] = MEM[5606] + MEM[9827];
assign MEM[13162] = MEM[5613] + MEM[6179];
assign MEM[13163] = MEM[5615] + MEM[7738];
assign MEM[13164] = MEM[5622] + MEM[7175];
assign MEM[13165] = MEM[5635] + MEM[3366];
assign MEM[13166] = MEM[5638] + MEM[6220];
assign MEM[13167] = MEM[5655] + MEM[7421];
assign MEM[13168] = MEM[5674] + MEM[8310];
assign MEM[13169] = MEM[5679] + MEM[9179];
assign MEM[13170] = MEM[5686] + MEM[3062];
assign MEM[13171] = MEM[5690] + MEM[876];
assign MEM[13172] = MEM[5694] + MEM[5702];
assign MEM[13173] = MEM[5700] + MEM[9065];
assign MEM[13174] = MEM[5707] + MEM[9042];
assign MEM[13175] = MEM[5711] + MEM[6404];
assign MEM[13176] = MEM[5715] + MEM[6484];
assign MEM[13177] = MEM[5732] + MEM[7343];
assign MEM[13178] = MEM[5733] + MEM[6173];
assign MEM[13179] = MEM[5734] + MEM[8822];
assign MEM[13180] = MEM[5735] + MEM[9102];
assign MEM[13181] = MEM[5742] + MEM[10762];
assign MEM[13182] = MEM[5749] + MEM[5210];
assign MEM[13183] = MEM[5751] + MEM[8303];
assign MEM[13184] = MEM[5757] + MEM[6692];
assign MEM[13185] = MEM[5759] + MEM[7213];
assign MEM[13186] = MEM[5762] + MEM[8564];
assign MEM[13187] = MEM[5765] + MEM[6999];
assign MEM[13188] = MEM[5770] + MEM[779];
assign MEM[13189] = MEM[5773] + MEM[11208];
assign MEM[13190] = MEM[5774] + MEM[9777];
assign MEM[13191] = MEM[5778] + MEM[6659];
assign MEM[13192] = MEM[5782] + MEM[6125];
assign MEM[13193] = MEM[5790] + MEM[6858];
assign MEM[13194] = MEM[5814] + MEM[7387];
assign MEM[13195] = MEM[5823] + MEM[8535];
assign MEM[13196] = MEM[5830] + MEM[2426];
assign MEM[13197] = MEM[5838] + MEM[7886];
assign MEM[13198] = MEM[5845] + MEM[4507];
assign MEM[13199] = MEM[5855] + MEM[9898];
assign MEM[13200] = MEM[5858] + MEM[10826];
assign MEM[13201] = MEM[5867] + MEM[7392];
assign MEM[13202] = MEM[5869] + MEM[10796];
assign MEM[13203] = MEM[5871] + MEM[7826];
assign MEM[13204] = MEM[5874] + MEM[10727];
assign MEM[13205] = MEM[5898] + MEM[6318];
assign MEM[13206] = MEM[5903] + MEM[10721];
assign MEM[13207] = MEM[5904] + MEM[10981];
assign MEM[13208] = MEM[5908] + MEM[7632];
assign MEM[13209] = MEM[5916] + MEM[2213];
assign MEM[13210] = MEM[5923] + MEM[8331];
assign MEM[13211] = MEM[5928] + MEM[6205];
assign MEM[13212] = MEM[5931] + MEM[5974];
assign MEM[13213] = MEM[5932] + MEM[7959];
assign MEM[13214] = MEM[5935] + MEM[6328];
assign MEM[13215] = MEM[5938] + MEM[10190];
assign MEM[13216] = MEM[5939] + MEM[7063];
assign MEM[13217] = MEM[5940] + MEM[7621];
assign MEM[13218] = MEM[5941] + MEM[782];
assign MEM[13219] = MEM[5950] + MEM[8040];
assign MEM[13220] = MEM[5951] + MEM[1879];
assign MEM[13221] = MEM[5956] + MEM[4962];
assign MEM[13222] = MEM[5964] + MEM[3807];
assign MEM[13223] = MEM[5966] + MEM[10712];
assign MEM[13224] = MEM[5967] + MEM[6859];
assign MEM[13225] = MEM[5970] + MEM[7717];
assign MEM[13226] = MEM[5972] + MEM[9588];
assign MEM[13227] = MEM[5979] + MEM[1275];
assign MEM[13228] = MEM[5980] + MEM[7767];
assign MEM[13229] = MEM[5990] + MEM[10373];
assign MEM[13230] = MEM[6005] + MEM[8819];
assign MEM[13231] = MEM[6012] + MEM[7218];
assign MEM[13232] = MEM[6015] + MEM[7504];
assign MEM[13233] = MEM[6021] + MEM[8245];
assign MEM[13234] = MEM[6023] + MEM[2483];
assign MEM[13235] = MEM[6045] + MEM[8174];
assign MEM[13236] = MEM[6055] + MEM[8537];
assign MEM[13237] = MEM[6087] + MEM[9181];
assign MEM[13238] = MEM[6093] + MEM[8828];
assign MEM[13239] = MEM[6094] + MEM[7244];
assign MEM[13240] = MEM[6103] + MEM[6795];
assign MEM[13241] = MEM[6107] + MEM[4077];
assign MEM[13242] = MEM[6131] + MEM[6481];
assign MEM[13243] = MEM[6132] + MEM[1639];
assign MEM[13244] = MEM[6143] + MEM[7999];
assign MEM[13245] = MEM[6158] + MEM[5982];
assign MEM[13246] = MEM[6159] + MEM[6360];
assign MEM[13247] = MEM[6164] + MEM[8339];
assign MEM[13248] = MEM[6165] + MEM[7754];
assign MEM[13249] = MEM[6171] + MEM[2524];
assign MEM[13250] = MEM[6178] + MEM[7235];
assign MEM[13251] = MEM[6191] + MEM[6246];
assign MEM[13252] = MEM[6195] + MEM[6744];
assign MEM[13253] = MEM[6196] + MEM[10656];
assign MEM[13254] = MEM[6198] + MEM[7076];
assign MEM[13255] = MEM[6199] + MEM[7084];
assign MEM[13256] = MEM[6211] + MEM[9324];
assign MEM[13257] = MEM[6214] + MEM[3636];
assign MEM[13258] = MEM[6221] + MEM[8455];
assign MEM[13259] = MEM[6227] + MEM[2311];
assign MEM[13260] = MEM[6231] + MEM[7873];
assign MEM[13261] = MEM[6237] + MEM[7734];
assign MEM[13262] = MEM[6238] + MEM[1227];
assign MEM[13263] = MEM[6239] + MEM[2559];
assign MEM[13264] = MEM[6254] + MEM[6957];
assign MEM[13265] = MEM[6261] + MEM[5991];
assign MEM[13266] = MEM[6263] + MEM[2188];
assign MEM[13267] = MEM[6272] + MEM[7167];
assign MEM[13268] = MEM[6275] + MEM[4535];
assign MEM[13269] = MEM[6282] + MEM[10578];
assign MEM[13270] = MEM[6307] + MEM[1027];
assign MEM[13271] = MEM[6309] + MEM[6391];
assign MEM[13272] = MEM[6313] + MEM[7344];
assign MEM[13273] = MEM[6332] + MEM[6985];
assign MEM[13274] = MEM[6336] + MEM[4146];
assign MEM[13275] = MEM[6342] + MEM[8270];
assign MEM[13276] = MEM[6346] + MEM[7898];
assign MEM[13277] = MEM[6347] + MEM[10621];
assign MEM[13278] = MEM[6348] + MEM[5650];
assign MEM[13279] = MEM[6361] + MEM[5798];
assign MEM[13280] = MEM[6365] + MEM[6814];
assign MEM[13281] = MEM[6371] + MEM[8087];
assign MEM[13282] = MEM[6379] + MEM[8622];
assign MEM[13283] = MEM[6388] + MEM[9388];
assign MEM[13284] = MEM[6409] + MEM[7144];
assign MEM[13285] = MEM[6411] + MEM[5174];
assign MEM[13286] = MEM[6414] + MEM[6694];
assign MEM[13287] = MEM[6415] + MEM[6556];
assign MEM[13288] = MEM[6424] + MEM[6463];
assign MEM[13289] = MEM[6443] + MEM[1676];
assign MEM[13290] = MEM[6445] + MEM[3019];
assign MEM[13291] = MEM[6462] + MEM[150];
assign MEM[13292] = MEM[6476] + MEM[10717];
assign MEM[13293] = MEM[6480] + MEM[7423];
assign MEM[13294] = MEM[6487] + MEM[11039];
assign MEM[13295] = MEM[6489] + MEM[7998];
assign MEM[13296] = MEM[6494] + MEM[8082];
assign MEM[13297] = MEM[6495] + MEM[7611];
assign MEM[13298] = MEM[6498] + MEM[10846];
assign MEM[13299] = MEM[6500] + MEM[7938];
assign MEM[13300] = MEM[6507] + MEM[7759];
assign MEM[13301] = MEM[6512] + MEM[10642];
assign MEM[13302] = MEM[6513] + MEM[1590];
assign MEM[13303] = MEM[6524] + MEM[4124];
assign MEM[13304] = MEM[6525] + MEM[10720];
assign MEM[13305] = MEM[6534] + MEM[6649];
assign MEM[13306] = MEM[6545] + MEM[8070];
assign MEM[13307] = MEM[6563] + MEM[7292];
assign MEM[13308] = MEM[6576] + MEM[6589];
assign MEM[13309] = MEM[6587] + MEM[4170];
assign MEM[13310] = MEM[6590] + MEM[9276];
assign MEM[13311] = MEM[6591] + MEM[10714];
assign MEM[13312] = MEM[6615] + MEM[2828];
assign MEM[13313] = MEM[6616] + MEM[8272];
assign MEM[13314] = MEM[6633] + MEM[2106];
assign MEM[13315] = MEM[6661] + MEM[948];
assign MEM[13316] = MEM[6669] + MEM[7248];
assign MEM[13317] = MEM[6671] + MEM[9814];
assign MEM[13318] = MEM[6677] + MEM[6969];
assign MEM[13319] = MEM[6686] + MEM[7345];
assign MEM[13320] = MEM[6691] + MEM[4515];
assign MEM[13321] = MEM[6700] + MEM[2067];
assign MEM[13322] = MEM[6701] + MEM[6808];
assign MEM[13323] = MEM[6708] + MEM[780];
assign MEM[13324] = MEM[6709] + MEM[1855];
assign MEM[13325] = MEM[6714] + MEM[7105];
assign MEM[13326] = MEM[6717] + MEM[3758];
assign MEM[13327] = MEM[6747] + MEM[2965];
assign MEM[13328] = MEM[6748] + MEM[9207];
assign MEM[13329] = MEM[6749] + MEM[2222];
assign MEM[13330] = MEM[6751] + MEM[6039];
assign MEM[13331] = MEM[6752] + MEM[8788];
assign MEM[13332] = MEM[6779] + MEM[8823];
assign MEM[13333] = MEM[6785] + MEM[6897];
assign MEM[13334] = MEM[6787] + MEM[7032];
assign MEM[13335] = MEM[6805] + MEM[1277];
assign MEM[13336] = MEM[6807] + MEM[8056];
assign MEM[13337] = MEM[6813] + MEM[4250];
assign MEM[13338] = MEM[6816] + MEM[7018];
assign MEM[13339] = MEM[6819] + MEM[7501];
assign MEM[13340] = MEM[6823] + MEM[7001];
assign MEM[13341] = MEM[6828] + MEM[8747];
assign MEM[13342] = MEM[6838] + MEM[3631];
assign MEM[13343] = MEM[6841] + MEM[7901];
assign MEM[13344] = MEM[6842] + MEM[7337];
assign MEM[13345] = MEM[6845] + MEM[6190];
assign MEM[13346] = MEM[6872] + MEM[7764];
assign MEM[13347] = MEM[6875] + MEM[8853];
assign MEM[13348] = MEM[6880] + MEM[8818];
assign MEM[13349] = MEM[6881] + MEM[7317];
assign MEM[13350] = MEM[6886] + MEM[8077];
assign MEM[13351] = MEM[6898] + MEM[7512];
assign MEM[13352] = MEM[6900] + MEM[8454];
assign MEM[13353] = MEM[6902] + MEM[4021];
assign MEM[13354] = MEM[6904] + MEM[10837];
assign MEM[13355] = MEM[6905] + MEM[7171];
assign MEM[13356] = MEM[6906] + MEM[10759];
assign MEM[13357] = MEM[6914] + MEM[10462];
assign MEM[13358] = MEM[6916] + MEM[6922];
assign MEM[13359] = MEM[6930] + MEM[7502];
assign MEM[13360] = MEM[6938] + MEM[8169];
assign MEM[13361] = MEM[6948] + MEM[10600];
assign MEM[13362] = MEM[6949] + MEM[335];
assign MEM[13363] = MEM[6951] + MEM[9264];
assign MEM[13364] = MEM[6958] + MEM[9191];
assign MEM[13365] = MEM[6959] + MEM[10735];
assign MEM[13366] = MEM[6964] + MEM[1031];
assign MEM[13367] = MEM[6968] + MEM[7622];
assign MEM[13368] = MEM[6970] + MEM[8870];
assign MEM[13369] = MEM[6972] + MEM[10728];
assign MEM[13370] = MEM[6980] + MEM[7295];
assign MEM[13371] = MEM[7004] + MEM[7279];
assign MEM[13372] = MEM[7024] + MEM[6212];
assign MEM[13373] = MEM[7027] + MEM[4138];
assign MEM[13374] = MEM[7031] + MEM[7737];
assign MEM[13375] = MEM[7036] + MEM[7885];
assign MEM[13376] = MEM[7040] + MEM[6353];
assign MEM[13377] = MEM[7047] + MEM[69];
assign MEM[13378] = MEM[7048] + MEM[8764];
assign MEM[13379] = MEM[7050] + MEM[4090];
assign MEM[13380] = MEM[7052] + MEM[2646];
assign MEM[13381] = MEM[7055] + MEM[6303];
assign MEM[13382] = MEM[7060] + MEM[6053];
assign MEM[13383] = MEM[7062] + MEM[7212];
assign MEM[13384] = MEM[7075] + MEM[5877];
assign MEM[13385] = MEM[7087] + MEM[8142];
assign MEM[13386] = MEM[7090] + MEM[867];
assign MEM[13387] = MEM[7112] + MEM[10028];
assign MEM[13388] = MEM[7124] + MEM[7732];
assign MEM[13389] = MEM[7132] + MEM[9948];
assign MEM[13390] = MEM[7134] + MEM[8043];
assign MEM[13391] = MEM[7138] + MEM[8757];
assign MEM[13392] = MEM[7142] + MEM[1844];
assign MEM[13393] = MEM[7147] + MEM[9182];
assign MEM[13394] = MEM[7149] + MEM[8559];
assign MEM[13395] = MEM[7161] + MEM[10056];
assign MEM[13396] = MEM[7166] + MEM[9806];
assign MEM[13397] = MEM[7179] + MEM[7306];
assign MEM[13398] = MEM[7198] + MEM[595];
assign MEM[13399] = MEM[7199] + MEM[7214];
assign MEM[13400] = MEM[7205] + MEM[7224];
assign MEM[13401] = MEM[7208] + MEM[2659];
assign MEM[13402] = MEM[7210] + MEM[7569];
assign MEM[13403] = MEM[7240] + MEM[8027];
assign MEM[13404] = MEM[7241] + MEM[8543];
assign MEM[13405] = MEM[7243] + MEM[2829];
assign MEM[13406] = MEM[7247] + MEM[8292];
assign MEM[13407] = MEM[7269] + MEM[7485];
assign MEM[13408] = MEM[7276] + MEM[8799];
assign MEM[13409] = MEM[7278] + MEM[6412];
assign MEM[13410] = MEM[7287] + MEM[8443];
assign MEM[13411] = MEM[7289] + MEM[8172];
assign MEM[13412] = MEM[7293] + MEM[7806];
assign MEM[13413] = MEM[7300] + MEM[563];
assign MEM[13414] = MEM[7301] + MEM[7602];
assign MEM[13415] = MEM[7302] + MEM[9739];
assign MEM[13416] = MEM[7304] + MEM[7757];
assign MEM[13417] = MEM[7307] + MEM[116];
assign MEM[13418] = MEM[7308] + MEM[3285];
assign MEM[13419] = MEM[7314] + MEM[5726];
assign MEM[13420] = MEM[7316] + MEM[4570];
assign MEM[13421] = MEM[7321] + MEM[9159];
assign MEM[13422] = MEM[7324] + MEM[9532];
assign MEM[13423] = MEM[7329] + MEM[10836];
assign MEM[13424] = MEM[7335] + MEM[9701];
assign MEM[13425] = MEM[7377] + MEM[7593];
assign MEM[13426] = MEM[7378] + MEM[7443];
assign MEM[13427] = MEM[7386] + MEM[1525];
assign MEM[13428] = MEM[7390] + MEM[6163];
assign MEM[13429] = MEM[7391] + MEM[7654];
assign MEM[13430] = MEM[7393] + MEM[7663];
assign MEM[13431] = MEM[7399] + MEM[8563];
assign MEM[13432] = MEM[7411] + MEM[3046];
assign MEM[13433] = MEM[7418] + MEM[6854];
assign MEM[13434] = MEM[7432] + MEM[7867];
assign MEM[13435] = MEM[7433] + MEM[7942];
assign MEM[13436] = MEM[7435] + MEM[9684];
assign MEM[13437] = MEM[7438] + MEM[11120];
assign MEM[13438] = MEM[7439] + MEM[8073];
assign MEM[13439] = MEM[7450] + MEM[7023];
assign MEM[13440] = MEM[7453] + MEM[10577];
assign MEM[13441] = MEM[7461] + MEM[94];
assign MEM[13442] = MEM[7463] + MEM[7594];
assign MEM[13443] = MEM[7469] + MEM[8201];
assign MEM[13444] = MEM[7476] + MEM[1203];
assign MEM[13445] = MEM[7484] + MEM[10752];
assign MEM[13446] = MEM[7490] + MEM[7596];
assign MEM[13447] = MEM[7507] + MEM[3543];
assign MEM[13448] = MEM[7517] + MEM[7892];
assign MEM[13449] = MEM[7522] + MEM[6312];
assign MEM[13450] = MEM[7529] + MEM[326];
assign MEM[13451] = MEM[7538] + MEM[7006];
assign MEM[13452] = MEM[7567] + MEM[10649];
assign MEM[13453] = MEM[7570] + MEM[2094];
assign MEM[13454] = MEM[7571] + MEM[7628];
assign MEM[13455] = MEM[7597] + MEM[7661];
assign MEM[13456] = MEM[7600] + MEM[10672];
assign MEM[13457] = MEM[7620] + MEM[8933];
assign MEM[13458] = MEM[7625] + MEM[10710];
assign MEM[13459] = MEM[7630] + MEM[8235];
assign MEM[13460] = MEM[7631] + MEM[10791];
assign MEM[13461] = MEM[7644] + MEM[6827];
assign MEM[13462] = MEM[7649] + MEM[8736];
assign MEM[13463] = MEM[7652] + MEM[8357];
assign MEM[13464] = MEM[7653] + MEM[8364];
assign MEM[13465] = MEM[7659] + MEM[7951];
assign MEM[13466] = MEM[7664] + MEM[7758];
assign MEM[13467] = MEM[7669] + MEM[5324];
assign MEM[13468] = MEM[7674] + MEM[6004];
assign MEM[13469] = MEM[7681] + MEM[5495];
assign MEM[13470] = MEM[7689] + MEM[3455];
assign MEM[13471] = MEM[7700] + MEM[3815];
assign MEM[13472] = MEM[7703] + MEM[2463];
assign MEM[13473] = MEM[7705] + MEM[4278];
assign MEM[13474] = MEM[7710] + MEM[10658];
assign MEM[13475] = MEM[7714] + MEM[9117];
assign MEM[13476] = MEM[7715] + MEM[4861];
assign MEM[13477] = MEM[7720] + MEM[1051];
assign MEM[13478] = MEM[7724] + MEM[4198];
assign MEM[13479] = MEM[7728] + MEM[8459];
assign MEM[13480] = MEM[7755] + MEM[2034];
assign MEM[13481] = MEM[7766] + MEM[6308];
assign MEM[13482] = MEM[7772] + MEM[4543];
assign MEM[13483] = MEM[7779] + MEM[7671];
assign MEM[13484] = MEM[7781] + MEM[7958];
assign MEM[13485] = MEM[7783] + MEM[4982];
assign MEM[13486] = MEM[7788] + MEM[8180];
assign MEM[13487] = MEM[7792] + MEM[9567];
assign MEM[13488] = MEM[7796] + MEM[6071];
assign MEM[13489] = MEM[7799] + MEM[10708];
assign MEM[13490] = MEM[7809] + MEM[8369];
assign MEM[13491] = MEM[7812] + MEM[8934];
assign MEM[13492] = MEM[7825] + MEM[7037];
assign MEM[13493] = MEM[7844] + MEM[5237];
assign MEM[13494] = MEM[7845] + MEM[10938];
assign MEM[13495] = MEM[7861] + MEM[10750];
assign MEM[13496] = MEM[7863] + MEM[10010];
assign MEM[13497] = MEM[7868] + MEM[4151];
assign MEM[13498] = MEM[7874] + MEM[7950];
assign MEM[13499] = MEM[7877] + MEM[9290];
assign MEM[13500] = MEM[7878] + MEM[8524];
assign MEM[13501] = MEM[7879] + MEM[7984];
assign MEM[13502] = MEM[7880] + MEM[1316];
assign MEM[13503] = MEM[7903] + MEM[9107];
assign MEM[13504] = MEM[7925] + MEM[5180];
assign MEM[13505] = MEM[7929] + MEM[10228];
assign MEM[13506] = MEM[7939] + MEM[9593];
assign MEM[13507] = MEM[7969] + MEM[2290];
assign MEM[13508] = MEM[7972] + MEM[167];
assign MEM[13509] = MEM[7981] + MEM[10998];
assign MEM[13510] = MEM[7987] + MEM[9043];
assign MEM[13511] = MEM[7988] + MEM[5930];
assign MEM[13512] = MEM[7992] + MEM[8221];
assign MEM[13513] = MEM[7997] + MEM[10693];
assign MEM[13514] = MEM[8003] + MEM[8987];
assign MEM[13515] = MEM[8008] + MEM[9426];
assign MEM[13516] = MEM[8013] + MEM[9148];
assign MEM[13517] = MEM[8019] + MEM[8243];
assign MEM[13518] = MEM[8020] + MEM[5710];
assign MEM[13519] = MEM[8021] + MEM[8253];
assign MEM[13520] = MEM[8025] + MEM[8740];
assign MEM[13521] = MEM[8034] + MEM[3907];
assign MEM[13522] = MEM[8050] + MEM[9157];
assign MEM[13523] = MEM[8053] + MEM[1780];
assign MEM[13524] = MEM[8054] + MEM[8640];
assign MEM[13525] = MEM[8062] + MEM[10724];
assign MEM[13526] = MEM[8063] + MEM[10500];
assign MEM[13527] = MEM[8083] + MEM[6325];
assign MEM[13528] = MEM[8088] + MEM[5300];
assign MEM[13529] = MEM[8105] + MEM[9053];
assign MEM[13530] = MEM[8106] + MEM[8118];
assign MEM[13531] = MEM[8115] + MEM[998];
assign MEM[13532] = MEM[8126] + MEM[7120];
assign MEM[13533] = MEM[8128] + MEM[5222];
assign MEM[13534] = MEM[8137] + MEM[8320];
assign MEM[13535] = MEM[8165] + MEM[6995];
assign MEM[13536] = MEM[8167] + MEM[8496];
assign MEM[13537] = MEM[8168] + MEM[9888];
assign MEM[13538] = MEM[8202] + MEM[5083];
assign MEM[13539] = MEM[8203] + MEM[6636];
assign MEM[13540] = MEM[8211] + MEM[11043];
assign MEM[13541] = MEM[8220] + MEM[9523];
assign MEM[13542] = MEM[8227] + MEM[4958];
assign MEM[13543] = MEM[8237] + MEM[8561];
assign MEM[13544] = MEM[8242] + MEM[9109];
assign MEM[13545] = MEM[8246] + MEM[8024];
assign MEM[13546] = MEM[8247] + MEM[11122];
assign MEM[13547] = MEM[8251] + MEM[9771];
assign MEM[13548] = MEM[8257] + MEM[8665];
assign MEM[13549] = MEM[8259] + MEM[9902];
assign MEM[13550] = MEM[8264] + MEM[10565];
assign MEM[13551] = MEM[8265] + MEM[4827];
assign MEM[13552] = MEM[8266] + MEM[9723];
assign MEM[13553] = MEM[8282] + MEM[634];
assign MEM[13554] = MEM[8284] + MEM[10844];
assign MEM[13555] = MEM[8286] + MEM[10692];
assign MEM[13556] = MEM[8291] + MEM[9832];
assign MEM[13557] = MEM[8294] + MEM[3998];
assign MEM[13558] = MEM[8299] + MEM[9568];
assign MEM[13559] = MEM[8301] + MEM[9186];
assign MEM[13560] = MEM[8302] + MEM[3759];
assign MEM[13561] = MEM[8306] + MEM[9347];
assign MEM[13562] = MEM[8319] + MEM[638];
assign MEM[13563] = MEM[8322] + MEM[3714];
assign MEM[13564] = MEM[8324] + MEM[8362];
assign MEM[13565] = MEM[8326] + MEM[10603];
assign MEM[13566] = MEM[8338] + MEM[8721];
assign MEM[13567] = MEM[8344] + MEM[6204];
assign MEM[13568] = MEM[8348] + MEM[10723];
assign MEM[13569] = MEM[8351] + MEM[5503];
assign MEM[13570] = MEM[8352] + MEM[7470];
assign MEM[13571] = MEM[8353] + MEM[9161];
assign MEM[13572] = MEM[8355] + MEM[10970];
assign MEM[13573] = MEM[8358] + MEM[9368];
assign MEM[13574] = MEM[8366] + MEM[4373];
assign MEM[13575] = MEM[8370] + MEM[8616];
assign MEM[13576] = MEM[8387] + MEM[10770];
assign MEM[13577] = MEM[8404] + MEM[7909];
assign MEM[13578] = MEM[8408] + MEM[10801];
assign MEM[13579] = MEM[8414] + MEM[10358];
assign MEM[13580] = MEM[8417] + MEM[8430];
assign MEM[13581] = MEM[8435] + MEM[10838];
assign MEM[13582] = MEM[8450] + MEM[8300];
assign MEM[13583] = MEM[8468] + MEM[3397];
assign MEM[13584] = MEM[8471] + MEM[7839];
assign MEM[13585] = MEM[8480] + MEM[10811];
assign MEM[13586] = MEM[8481] + MEM[9145];
assign MEM[13587] = MEM[8500] + MEM[8536];
assign MEM[13588] = MEM[8516] + MEM[6135];
assign MEM[13589] = MEM[8519] + MEM[8287];
assign MEM[13590] = MEM[8521] + MEM[9285];
assign MEM[13591] = MEM[8538] + MEM[8445];
assign MEM[13592] = MEM[8553] + MEM[5771];
assign MEM[13593] = MEM[8572] + MEM[10627];
assign MEM[13594] = MEM[8582] + MEM[7038];
assign MEM[13595] = MEM[8620] + MEM[7607];
assign MEM[13596] = MEM[8639] + MEM[10487];
assign MEM[13597] = MEM[8662] + MEM[10645];
assign MEM[13598] = MEM[8663] + MEM[5859];
assign MEM[13599] = MEM[8666] + MEM[7937];
assign MEM[13600] = MEM[8679] + MEM[10726];
assign MEM[13601] = MEM[8681] + MEM[4453];
assign MEM[13602] = MEM[8683] + MEM[2475];
assign MEM[13603] = MEM[8685] + MEM[10911];
assign MEM[13604] = MEM[8688] + MEM[10843];
assign MEM[13605] = MEM[8689] + MEM[4315];
assign MEM[13606] = MEM[8697] + MEM[3775];
assign MEM[13607] = MEM[8705] + MEM[10559];
assign MEM[13608] = MEM[8716] + MEM[6285];
assign MEM[13609] = MEM[8722] + MEM[10715];
assign MEM[13610] = MEM[8724] + MEM[7900];
assign MEM[13611] = MEM[8726] + MEM[9672];
assign MEM[13612] = MEM[8730] + MEM[4358];
assign MEM[13613] = MEM[8731] + MEM[10531];
assign MEM[13614] = MEM[8758] + MEM[2230];
assign MEM[13615] = MEM[8761] + MEM[10876];
assign MEM[13616] = MEM[8777] + MEM[5383];
assign MEM[13617] = MEM[8784] + MEM[2494];
assign MEM[13618] = MEM[8798] + MEM[9995];
assign MEM[13619] = MEM[8832] + MEM[10659];
assign MEM[13620] = MEM[8837] + MEM[9835];
assign MEM[13621] = MEM[8838] + MEM[3887];
assign MEM[13622] = MEM[8857] + MEM[3934];
assign MEM[13623] = MEM[8879] + MEM[7191];
assign MEM[13624] = MEM[8883] + MEM[8807];
assign MEM[13625] = MEM[8912] + MEM[10608];
assign MEM[13626] = MEM[8923] + MEM[7760];
assign MEM[13627] = MEM[8928] + MEM[7338];
assign MEM[13628] = MEM[8930] + MEM[9728];
assign MEM[13629] = MEM[8937] + MEM[615];
assign MEM[13630] = MEM[8951] + MEM[7176];
assign MEM[13631] = MEM[8954] + MEM[8055];
assign MEM[13632] = MEM[8974] + MEM[197];
assign MEM[13633] = MEM[8991] + MEM[2645];
assign MEM[13634] = MEM[9007] + MEM[6115];
assign MEM[13635] = MEM[9018] + MEM[9188];
assign MEM[13636] = MEM[9077] + MEM[10733];
assign MEM[13637] = MEM[9086] + MEM[10530];
assign MEM[13638] = MEM[9091] + MEM[10855];
assign MEM[13639] = MEM[9094] + MEM[7655];
assign MEM[13640] = MEM[9127] + MEM[6743];
assign MEM[13641] = MEM[9137] + MEM[8796];
assign MEM[13642] = MEM[9149] + MEM[262];
assign MEM[13643] = MEM[9184] + MEM[4775];
assign MEM[13644] = MEM[9204] + MEM[4054];
assign MEM[13645] = MEM[9228] + MEM[9648];
assign MEM[13646] = MEM[9229] + MEM[9706];
assign MEM[13647] = MEM[9247] + MEM[10797];
assign MEM[13648] = MEM[9265] + MEM[10691];
assign MEM[13649] = MEM[9280] + MEM[4047];
assign MEM[13650] = MEM[9286] + MEM[8596];
assign MEM[13651] = MEM[9306] + MEM[10858];
assign MEM[13652] = MEM[9353] + MEM[2252];
assign MEM[13653] = MEM[9371] + MEM[918];
assign MEM[13654] = MEM[9378] + MEM[8273];
assign MEM[13655] = MEM[9389] + MEM[8738];
assign MEM[13656] = MEM[9419] + MEM[2958];
assign MEM[13657] = MEM[9453] + MEM[8829];
assign MEM[13658] = MEM[9494] + MEM[5142];
assign MEM[13659] = MEM[9507] + MEM[7773];
assign MEM[13660] = MEM[9531] + MEM[9309];
assign MEM[13661] = MEM[9537] + MEM[10809];
assign MEM[13662] = MEM[9543] + MEM[10624];
assign MEM[13663] = MEM[9549] + MEM[4765];
assign MEM[13664] = MEM[9570] + MEM[4180];
assign MEM[13665] = MEM[9585] + MEM[10973];
assign MEM[13666] = MEM[9591] + MEM[10833];
assign MEM[13667] = MEM[9604] + MEM[2459];
assign MEM[13668] = MEM[9612] + MEM[10780];
assign MEM[13669] = MEM[9616] + MEM[9743];
assign MEM[13670] = MEM[9625] + MEM[10793];
assign MEM[13671] = MEM[9650] + MEM[7496];
assign MEM[13672] = MEM[9652] + MEM[7716];
assign MEM[13673] = MEM[9659] + MEM[3365];
assign MEM[13674] = MEM[9676] + MEM[6982];
assign MEM[13675] = MEM[9709] + MEM[11263];
assign MEM[13676] = MEM[9753] + MEM[10897];
assign MEM[13677] = MEM[9769] + MEM[10831];
assign MEM[13678] = MEM[9788] + MEM[10862];
assign MEM[13679] = MEM[9980] + MEM[10881];
assign MEM[13680] = MEM[10134] + MEM[5662];
assign MEM[13681] = MEM[10569] + MEM[5654];
assign MEM[13682] = MEM[10574] + MEM[8675];
assign MEM[13683] = MEM[10575] + MEM[9998];
assign MEM[13684] = MEM[10576] + MEM[7546];
assign MEM[13685] = MEM[10593] + MEM[7846];
assign MEM[13686] = MEM[10595] + MEM[10220];
assign MEM[13687] = MEM[10602] + MEM[4786];
assign MEM[13688] = MEM[10607] + MEM[389];
assign MEM[13689] = MEM[10619] + MEM[7088];
assign MEM[13690] = MEM[10623] + MEM[1394];
assign MEM[13691] = MEM[10633] + MEM[7798];
assign MEM[13692] = MEM[10644] + MEM[988];
assign MEM[13693] = MEM[10664] + MEM[8759];
assign MEM[13694] = MEM[10671] + MEM[55];
assign MEM[13695] = MEM[10674] + MEM[9433];
assign MEM[13696] = MEM[10681] + MEM[453];
assign MEM[13697] = MEM[10682] + MEM[5839];
assign MEM[13698] = MEM[10688] + MEM[5070];
assign MEM[13699] = MEM[10694] + MEM[2006];
assign MEM[13700] = MEM[10699] + MEM[10192];
assign MEM[13701] = MEM[10737] + MEM[3165];
assign MEM[13702] = MEM[10738] + MEM[6491];
assign MEM[13703] = MEM[10739] + MEM[1047];
assign MEM[13704] = MEM[10743] + MEM[2686];
assign MEM[13705] = MEM[10744] + MEM[1730];
assign MEM[13706] = MEM[10745] + MEM[9505];
assign MEM[13707] = MEM[10746] + MEM[10971];
assign MEM[13708] = MEM[10747] + MEM[2047];
assign MEM[13709] = MEM[10748] + MEM[3788];
assign MEM[13710] = MEM[10753] + MEM[1994];
assign MEM[13711] = MEM[10755] + MEM[2557];
assign MEM[13712] = MEM[10756] + MEM[78];
assign MEM[13713] = MEM[10757] + MEM[8413];
assign MEM[13714] = MEM[10763] + MEM[7100];
assign MEM[13715] = MEM[10765] + MEM[1757];
assign MEM[13716] = MEM[10769] + MEM[8065];
assign MEM[13717] = MEM[10774] + MEM[7054];
assign MEM[13718] = MEM[10775] + MEM[10840];
assign MEM[13719] = MEM[10778] + MEM[5271];
assign MEM[13720] = MEM[10779] + MEM[11251];
assign MEM[13721] = MEM[10781] + MEM[6492];
assign MEM[13722] = MEM[10782] + MEM[223];
assign MEM[13723] = MEM[10784] + MEM[5043];
assign MEM[13724] = MEM[10786] + MEM[10143];
assign MEM[13725] = MEM[10792] + MEM[1147];
assign MEM[13726] = MEM[10798] + MEM[3530];
assign MEM[13727] = MEM[10800] + MEM[8173];
assign MEM[13728] = MEM[10802] + MEM[5772];
assign MEM[13729] = MEM[10803] + MEM[5630];
assign MEM[13730] = MEM[10804] + MEM[1940];
assign MEM[13731] = MEM[10805] + MEM[794];
assign MEM[13732] = MEM[10807] + MEM[1645];
assign MEM[13733] = MEM[10814] + MEM[2717];
assign MEM[13734] = MEM[10815] + MEM[1234];
assign MEM[13735] = MEM[10816] + MEM[10829];
assign MEM[13736] = MEM[10818] + MEM[2205];
assign MEM[13737] = MEM[10819] + MEM[5022];
assign MEM[13738] = MEM[10821] + MEM[5100];
assign MEM[13739] = MEM[10823] + MEM[3012];
assign MEM[13740] = MEM[10825] + MEM[4661];
assign MEM[13741] = MEM[10828] + MEM[8545];
assign MEM[13742] = MEM[10830] + MEM[9327];
assign MEM[13743] = MEM[10842] + MEM[869];
assign MEM[13744] = MEM[10845] + MEM[8577];
assign MEM[13745] = MEM[10847] + MEM[8120];
assign MEM[13746] = MEM[10848] + MEM[7310];
assign MEM[13747] = MEM[10851] + MEM[9062];
assign MEM[13748] = MEM[10852] + MEM[7530];
assign MEM[13749] = MEM[10854] + MEM[7058];
assign MEM[13750] = MEM[10857] + MEM[8748];
assign MEM[13751] = MEM[10860] + MEM[8978];
assign MEM[13752] = MEM[10867] + MEM[3926];
assign MEM[13753] = MEM[10868] + MEM[2347];
assign MEM[13754] = MEM[10869] + MEM[5339];
assign MEM[13755] = MEM[10870] + MEM[7578];
assign MEM[13756] = MEM[10871] + MEM[6652];
assign MEM[13757] = MEM[10872] + MEM[2940];
assign MEM[13758] = MEM[10873] + MEM[11023];
assign MEM[13759] = MEM[10875] + MEM[629];
assign MEM[13760] = MEM[10884] + MEM[788];
assign MEM[13761] = MEM[10885] + MEM[7366];
assign MEM[13762] = MEM[10886] + MEM[4405];
assign MEM[13763] = MEM[10887] + MEM[7794];
assign MEM[13764] = MEM[10891] + MEM[8097];
assign MEM[13765] = MEM[10893] + MEM[7242];
assign MEM[13766] = MEM[10895] + MEM[7971];
assign MEM[13767] = MEM[10899] + MEM[1279];
assign MEM[13768] = MEM[10902] + MEM[5983];
assign MEM[13769] = MEM[10904] + MEM[10935];
assign MEM[13770] = MEM[10905] + MEM[2711];
assign MEM[13771] = MEM[10908] + MEM[2547];
assign MEM[13772] = MEM[10910] + MEM[8359];
assign MEM[13773] = MEM[10917] + MEM[8506];
assign MEM[13774] = MEM[10918] + MEM[8626];
assign MEM[13775] = MEM[10919] + MEM[575];
assign MEM[13776] = MEM[10922] + MEM[2194];
assign MEM[13777] = MEM[10934] + MEM[10309];
assign MEM[13778] = MEM[10936] + MEM[7606];
assign MEM[13779] = MEM[10937] + MEM[4710];
assign MEM[13780] = MEM[10946] + MEM[4252];
assign MEM[13781] = MEM[10947] + MEM[9506];
assign MEM[13782] = MEM[10948] + MEM[4171];
assign MEM[13783] = MEM[10950] + MEM[6293];
assign MEM[13784] = MEM[10956] + MEM[3532];
assign MEM[13785] = MEM[10959] + MEM[807];
assign MEM[13786] = MEM[10962] + MEM[8767];
assign MEM[13787] = MEM[10964] + MEM[5919];
assign MEM[13788] = MEM[10967] + MEM[7683];
assign MEM[13789] = MEM[10969] + MEM[2118];
assign MEM[13790] = MEM[10976] + MEM[9465];
assign MEM[13791] = MEM[10978] + MEM[6298];
assign MEM[13792] = MEM[10982] + MEM[8427];
assign MEM[13793] = MEM[10985] + MEM[1468];
assign MEM[13794] = MEM[10986] + MEM[7139];
assign MEM[13795] = MEM[10988] + MEM[11044];
assign MEM[13796] = MEM[10989] + MEM[2062];
assign MEM[13797] = MEM[10990] + MEM[1395];
assign MEM[13798] = MEM[10993] + MEM[7159];
assign MEM[13799] = MEM[10994] + MEM[10900];
assign MEM[13800] = MEM[10996] + MEM[10059];
assign MEM[13801] = MEM[11001] + MEM[9216];
assign MEM[13802] = MEM[11003] + MEM[9190];
assign MEM[13803] = MEM[11007] + MEM[5598];
assign MEM[13804] = MEM[11010] + MEM[7657];
assign MEM[13805] = MEM[11011] + MEM[542];
assign MEM[13806] = MEM[11012] + MEM[7456];
assign MEM[13807] = MEM[11017] + MEM[8233];
assign MEM[13808] = MEM[11018] + MEM[3918];
assign MEM[13809] = MEM[11022] + MEM[2925];
assign MEM[13810] = MEM[11025] + MEM[8171];
assign MEM[13811] = MEM[11026] + MEM[8032];
assign MEM[13812] = MEM[11030] + MEM[4517];
assign MEM[13813] = MEM[11068] + MEM[3738];
assign MEM[13814] = MEM[11081] + MEM[2173];
assign MEM[13815] = MEM[11086] + MEM[2119];
assign MEM[13816] = MEM[11097] + MEM[8772];
assign MEM[13817] = MEM[11099] + MEM[9113];
assign MEM[13818] = MEM[11104] + MEM[2579];
assign MEM[13819] = MEM[11108] + MEM[8067];
assign MEM[13820] = MEM[11116] + MEM[8739];
assign MEM[13821] = MEM[11131] + MEM[1022];
assign MEM[13822] = MEM[11155] + MEM[2631];
assign MEM[13823] = MEM[11169] + MEM[3404];
assign MEM[13824] = MEM[11184] + MEM[8398];
assign MEM[13825] = MEM[11290] + MEM[9060];
assign MEM[13826] = MEM[12847] + MEM[11239];
assign MEM[13827] = MEM[7] + MEM[8181];
assign MEM[13828] = MEM[38] + MEM[1861];
assign MEM[13829] = MEM[53] + MEM[3110];
assign MEM[13830] = MEM[54] + MEM[3874];
assign MEM[13831] = MEM[61] + MEM[903];
assign MEM[13832] = MEM[62] + MEM[8317];
assign MEM[13833] = MEM[63] + MEM[862];
assign MEM[13834] = MEM[71] + MEM[7840];
assign MEM[13835] = MEM[79] + MEM[3994];
assign MEM[13836] = MEM[93] + MEM[5786];
assign MEM[13837] = MEM[102] + MEM[4652];
assign MEM[13838] = MEM[103] + MEM[3844];
assign MEM[13839] = MEM[107] + MEM[350];
assign MEM[13840] = MEM[110] + MEM[1271];
assign MEM[13841] = MEM[157] + MEM[1331];
assign MEM[13842] = MEM[158] + MEM[2298];
assign MEM[13843] = MEM[181] + MEM[1724];
assign MEM[13844] = MEM[182] + MEM[1318];
assign MEM[13845] = MEM[191] + MEM[4388];
assign MEM[13846] = MEM[205] + MEM[8285];
assign MEM[13847] = MEM[206] + MEM[4123];
assign MEM[13848] = MEM[213] + MEM[342];
assign MEM[13849] = MEM[214] + MEM[2803];
assign MEM[13850] = MEM[229] + MEM[4549];
assign MEM[13851] = MEM[238] + MEM[7888];
assign MEM[13852] = MEM[246] + MEM[2860];
assign MEM[13853] = MEM[261] + MEM[5020];
assign MEM[13854] = MEM[270] + MEM[828];
assign MEM[13855] = MEM[278] + MEM[8297];
assign MEM[13856] = MEM[283] + MEM[11111];
assign MEM[13857] = MEM[285] + MEM[9581];
assign MEM[13858] = MEM[292] + MEM[2618];
assign MEM[13859] = MEM[300] + MEM[4222];
assign MEM[13860] = MEM[303] + MEM[2086];
assign MEM[13861] = MEM[319] + MEM[2599];
assign MEM[13862] = MEM[325] + MEM[1099];
assign MEM[13863] = MEM[327] + MEM[8586];
assign MEM[13864] = MEM[347] + MEM[7923];
assign MEM[13865] = MEM[348] + MEM[2446];
assign MEM[13866] = MEM[356] + MEM[4229];
assign MEM[13867] = MEM[362] + MEM[1725];
assign MEM[13868] = MEM[367] + MEM[3159];
assign MEM[13869] = MEM[374] + MEM[855];
assign MEM[13870] = MEM[379] + MEM[1222];
assign MEM[13871] = MEM[382] + MEM[1055];
assign MEM[13872] = MEM[388] + MEM[1614];
assign MEM[13873] = MEM[390] + MEM[4894];
assign MEM[13874] = MEM[390] + MEM[5087];
assign MEM[13875] = MEM[391] + MEM[7057];
assign MEM[13876] = MEM[397] + MEM[7353];
assign MEM[13877] = MEM[398] + MEM[10866];
assign MEM[13878] = MEM[403] + MEM[3747];
assign MEM[13879] = MEM[404] + MEM[5327];
assign MEM[13880] = MEM[411] + MEM[2215];
assign MEM[13881] = MEM[412] + MEM[2462];
assign MEM[13882] = MEM[413] + MEM[6380];
assign MEM[13883] = MEM[437] + MEM[2819];
assign MEM[13884] = MEM[439] + MEM[2811];
assign MEM[13885] = MEM[446] + MEM[3020];
assign MEM[13886] = MEM[461] + MEM[7904];
assign MEM[13887] = MEM[478] + MEM[3955];
assign MEM[13888] = MEM[485] + MEM[719];
assign MEM[13889] = MEM[486] + MEM[5470];
assign MEM[13890] = MEM[499] + MEM[8145];
assign MEM[13891] = MEM[502] + MEM[1582];
assign MEM[13892] = MEM[508] + MEM[1326];
assign MEM[13893] = MEM[510] + MEM[2870];
assign MEM[13894] = MEM[511] + MEM[3550];
assign MEM[13895] = MEM[535] + MEM[3173];
assign MEM[13896] = MEM[539] + MEM[7355];
assign MEM[13897] = MEM[557] + MEM[1558];
assign MEM[13898] = MEM[565] + MEM[7072];
assign MEM[13899] = MEM[567] + MEM[3223];
assign MEM[13900] = MEM[572] + MEM[3060];
assign MEM[13901] = MEM[578] + MEM[2059];
assign MEM[13902] = MEM[585] + MEM[6431];
assign MEM[13903] = MEM[587] + MEM[8135];
assign MEM[13904] = MEM[590] + MEM[8179];
assign MEM[13905] = MEM[599] + MEM[7074];
assign MEM[13906] = MEM[600] + MEM[7151];
assign MEM[13907] = MEM[601] + MEM[3325];
assign MEM[13908] = MEM[605] + MEM[1034];
assign MEM[13909] = MEM[606] + MEM[2814];
assign MEM[13910] = MEM[606] + MEM[11363];
assign MEM[13911] = MEM[612] + MEM[4805];
assign MEM[13912] = MEM[613] + MEM[5430];
assign MEM[13913] = MEM[619] + MEM[3188];
assign MEM[13914] = MEM[623] + MEM[7357];
assign MEM[13915] = MEM[630] + MEM[2078];
assign MEM[13916] = MEM[637] + MEM[979];
assign MEM[13917] = MEM[644] + MEM[1133];
assign MEM[13918] = MEM[645] + MEM[9361];
assign MEM[13919] = MEM[646] + MEM[748];
assign MEM[13920] = MEM[654] + MEM[4679];
assign MEM[13921] = MEM[662] + MEM[3876];
assign MEM[13922] = MEM[671] + MEM[3245];
assign MEM[13923] = MEM[679] + MEM[8651];
assign MEM[13924] = MEM[685] + MEM[3847];
assign MEM[13925] = MEM[686] + MEM[5030];
assign MEM[13926] = MEM[694] + MEM[5069];
assign MEM[13927] = MEM[701] + MEM[3878];
assign MEM[13928] = MEM[702] + MEM[826];
assign MEM[13929] = MEM[717] + MEM[7768];
assign MEM[13930] = MEM[718] + MEM[1228];
assign MEM[13931] = MEM[735] + MEM[7275];
assign MEM[13932] = MEM[739] + MEM[3315];
assign MEM[13933] = MEM[740] + MEM[5298];
assign MEM[13934] = MEM[745] + MEM[7678];
assign MEM[13935] = MEM[749] + MEM[3861];
assign MEM[13936] = MEM[750] + MEM[1931];
assign MEM[13937] = MEM[751] + MEM[1819];
assign MEM[13938] = MEM[757] + MEM[3351];
assign MEM[13939] = MEM[760] + MEM[7656];
assign MEM[13940] = MEM[763] + MEM[2795];
assign MEM[13941] = MEM[773] + MEM[3773];
assign MEM[13942] = MEM[778] + MEM[2787];
assign MEM[13943] = MEM[783] + MEM[9366];
assign MEM[13944] = MEM[786] + MEM[5807];
assign MEM[13945] = MEM[787] + MEM[4726];
assign MEM[13946] = MEM[791] + MEM[3199];
assign MEM[13947] = MEM[797] + MEM[3316];
assign MEM[13948] = MEM[798] + MEM[1045];
assign MEM[13949] = MEM[799] + MEM[2971];
assign MEM[13950] = MEM[802] + MEM[2789];
assign MEM[13951] = MEM[805] + MEM[3334];
assign MEM[13952] = MEM[815] + MEM[3619];
assign MEM[13953] = MEM[819] + MEM[2388];
assign MEM[13954] = MEM[829] + MEM[3326];
assign MEM[13955] = MEM[839] + MEM[2434];
assign MEM[13956] = MEM[842] + MEM[3412];
assign MEM[13957] = MEM[843] + MEM[6337];
assign MEM[13958] = MEM[844] + MEM[8170];
assign MEM[13959] = MEM[852] + MEM[4379];
assign MEM[13960] = MEM[868] + MEM[3910];
assign MEM[13961] = MEM[871] + MEM[3342];
assign MEM[13962] = MEM[874] + MEM[1766];
assign MEM[13963] = MEM[909] + MEM[7197];
assign MEM[13964] = MEM[916] + MEM[8762];
assign MEM[13965] = MEM[919] + MEM[5747];
assign MEM[13966] = MEM[926] + MEM[7572];
assign MEM[13967] = MEM[931] + MEM[3172];
assign MEM[13968] = MEM[933] + MEM[8692];
assign MEM[13969] = MEM[935] + MEM[4742];
assign MEM[13970] = MEM[938] + MEM[3735];
assign MEM[13971] = MEM[943] + MEM[11470];
assign MEM[13972] = MEM[951] + MEM[7982];
assign MEM[13973] = MEM[975] + MEM[1286];
assign MEM[13974] = MEM[995] + MEM[8615];
assign MEM[13975] = MEM[996] + MEM[3460];
assign MEM[13976] = MEM[1011] + MEM[4074];
assign MEM[13977] = MEM[1013] + MEM[1188];
assign MEM[13978] = MEM[1014] + MEM[3739];
assign MEM[13979] = MEM[1018] + MEM[2182];
assign MEM[13980] = MEM[1019] + MEM[8658];
assign MEM[13981] = MEM[1035] + MEM[5748];
assign MEM[13982] = MEM[1038] + MEM[6831];
assign MEM[13983] = MEM[1042] + MEM[2279];
assign MEM[13984] = MEM[1050] + MEM[2844];
assign MEM[13985] = MEM[1078] + MEM[7383];
assign MEM[13986] = MEM[1079] + MEM[8256];
assign MEM[13987] = MEM[1082] + MEM[6422];
assign MEM[13988] = MEM[1085] + MEM[7479];
assign MEM[13989] = MEM[1086] + MEM[9839];
assign MEM[13990] = MEM[1092] + MEM[5900];
assign MEM[13991] = MEM[1101] + MEM[7968];
assign MEM[13992] = MEM[1118] + MEM[1589];
assign MEM[13993] = MEM[1127] + MEM[9160];
assign MEM[13994] = MEM[1141] + MEM[1597];
assign MEM[13995] = MEM[1143] + MEM[6988];
assign MEM[13996] = MEM[1149] + MEM[7413];
assign MEM[13997] = MEM[1154] + MEM[4172];
assign MEM[13998] = MEM[1162] + MEM[1807];
assign MEM[13999] = MEM[1167] + MEM[9431];
assign MEM[14000] = MEM[1170] + MEM[7434];
assign MEM[14001] = MEM[1179] + MEM[10841];
assign MEM[14002] = MEM[1183] + MEM[2989];
assign MEM[14003] = MEM[1183] + MEM[8670];
assign MEM[14004] = MEM[1199] + MEM[2555];
assign MEM[14005] = MEM[1204] + MEM[2818];
assign MEM[14006] = MEM[1205] + MEM[8598];
assign MEM[14007] = MEM[1206] + MEM[10347];
assign MEM[14008] = MEM[1215] + MEM[7146];
assign MEM[14009] = MEM[1220] + MEM[5779];
assign MEM[14010] = MEM[1229] + MEM[7978];
assign MEM[14011] = MEM[1243] + MEM[9772];
assign MEM[14012] = MEM[1261] + MEM[5003];
assign MEM[14013] = MEM[1266] + MEM[5623];
assign MEM[14014] = MEM[1267] + MEM[1388];
assign MEM[14015] = MEM[1269] + MEM[7670];
assign MEM[14016] = MEM[1282] + MEM[4503];
assign MEM[14017] = MEM[1283] + MEM[7941];
assign MEM[14018] = MEM[1285] + MEM[1378];
assign MEM[14019] = MEM[1287] + MEM[3382];
assign MEM[14020] = MEM[1291] + MEM[4300];
assign MEM[14021] = MEM[1295] + MEM[2947];
assign MEM[14022] = MEM[1299] + MEM[8469];
assign MEM[14023] = MEM[1300] + MEM[8308];
assign MEM[14024] = MEM[1306] + MEM[1699];
assign MEM[14025] = MEM[1307] + MEM[1534];
assign MEM[14026] = MEM[1310] + MEM[6538];
assign MEM[14027] = MEM[1311] + MEM[1781];
assign MEM[14028] = MEM[1317] + MEM[2365];
assign MEM[14029] = MEM[1319] + MEM[1830];
assign MEM[14030] = MEM[1323] + MEM[2733];
assign MEM[14031] = MEM[1343] + MEM[4410];
assign MEM[14032] = MEM[1350] + MEM[3095];
assign MEM[14033] = MEM[1351] + MEM[7462];
assign MEM[14034] = MEM[1357] + MEM[5060];
assign MEM[14035] = MEM[1359] + MEM[5629];
assign MEM[14036] = MEM[1372] + MEM[4005];
assign MEM[14037] = MEM[1373] + MEM[6362];
assign MEM[14038] = MEM[1382] + MEM[7748];
assign MEM[14039] = MEM[1383] + MEM[1662];
assign MEM[14040] = MEM[1391] + MEM[3373];
assign MEM[14041] = MEM[1399] + MEM[2831];
assign MEM[14042] = MEM[1402] + MEM[3092];
assign MEM[14043] = MEM[1413] + MEM[6029];
assign MEM[14044] = MEM[1419] + MEM[5255];
assign MEM[14045] = MEM[1421] + MEM[2005];
assign MEM[14046] = MEM[1430] + MEM[4682];
assign MEM[14047] = MEM[1436] + MEM[7782];
assign MEM[14048] = MEM[1442] + MEM[8240];
assign MEM[14049] = MEM[1450] + MEM[3109];
assign MEM[14050] = MEM[1452] + MEM[8429];
assign MEM[14051] = MEM[1458] + MEM[1738];
assign MEM[14052] = MEM[1471] + MEM[2586];
assign MEM[14053] = MEM[1474] + MEM[9068];
assign MEM[14054] = MEM[1476] + MEM[3522];
assign MEM[14055] = MEM[1477] + MEM[5202];
assign MEM[14056] = MEM[1482] + MEM[6943];
assign MEM[14057] = MEM[1486] + MEM[3044];
assign MEM[14058] = MEM[1491] + MEM[9812];
assign MEM[14059] = MEM[1494] + MEM[9101];
assign MEM[14060] = MEM[1495] + MEM[2772];
assign MEM[14061] = MEM[1499] + MEM[10974];
assign MEM[14062] = MEM[1506] + MEM[2623];
assign MEM[14063] = MEM[1510] + MEM[5364];
assign MEM[14064] = MEM[1511] + MEM[6578];
assign MEM[14065] = MEM[1515] + MEM[4235];
assign MEM[14066] = MEM[1517] + MEM[7096];
assign MEM[14067] = MEM[1519] + MEM[6837];
assign MEM[14068] = MEM[1524] + MEM[2238];
assign MEM[14069] = MEM[1535] + MEM[6117];
assign MEM[14070] = MEM[1541] + MEM[1852];
assign MEM[14071] = MEM[1542] + MEM[5126];
assign MEM[14072] = MEM[1547] + MEM[3626];
assign MEM[14073] = MEM[1573] + MEM[6588];
assign MEM[14074] = MEM[1588] + MEM[8585];
assign MEM[14075] = MEM[1610] + MEM[2908];
assign MEM[14076] = MEM[1611] + MEM[5764];
assign MEM[14077] = MEM[1613] + MEM[7141];
assign MEM[14078] = MEM[1621] + MEM[6323];
assign MEM[14079] = MEM[1623] + MEM[2191];
assign MEM[14080] = MEM[1627] + MEM[7061];
assign MEM[14081] = MEM[1631] + MEM[3142];
assign MEM[14082] = MEM[1634] + MEM[4243];
assign MEM[14083] = MEM[1635] + MEM[4301];
assign MEM[14084] = MEM[1651] + MEM[11032];
assign MEM[14085] = MEM[1655] + MEM[9308];
assign MEM[14086] = MEM[1667] + MEM[2354];
assign MEM[14087] = MEM[1674] + MEM[5151];
assign MEM[14088] = MEM[1682] + MEM[10931];
assign MEM[14089] = MEM[1683] + MEM[4595];
assign MEM[14090] = MEM[1690] + MEM[5131];
assign MEM[14091] = MEM[1691] + MEM[3764];
assign MEM[14092] = MEM[1692] + MEM[9910];
assign MEM[14093] = MEM[1693] + MEM[3358];
assign MEM[14094] = MEM[1701] + MEM[2139];
assign MEM[14095] = MEM[1703] + MEM[5038];
assign MEM[14096] = MEM[1706] + MEM[3054];
assign MEM[14097] = MEM[1709] + MEM[2447];
assign MEM[14098] = MEM[1711] + MEM[4996];
assign MEM[14099] = MEM[1718] + MEM[4802];
assign MEM[14100] = MEM[1733] + MEM[2927];
assign MEM[14101] = MEM[1738] + MEM[7699];
assign MEM[14102] = MEM[1746] + MEM[2164];
assign MEM[14103] = MEM[1790] + MEM[5994];
assign MEM[14104] = MEM[1806] + MEM[1965];
assign MEM[14105] = MEM[1827] + MEM[9251];
assign MEM[14106] = MEM[1847] + MEM[4516];
assign MEM[14107] = MEM[1867] + MEM[8010];
assign MEM[14108] = MEM[1869] + MEM[2882];
assign MEM[14109] = MEM[1883] + MEM[2986];
assign MEM[14110] = MEM[1885] + MEM[9238];
assign MEM[14111] = MEM[1915] + MEM[7876];
assign MEM[14112] = MEM[1917] + MEM[6839];
assign MEM[14113] = MEM[1922] + MEM[10013];
assign MEM[14114] = MEM[1924] + MEM[2741];
assign MEM[14115] = MEM[1925] + MEM[5342];
assign MEM[14116] = MEM[1933] + MEM[2589];
assign MEM[14117] = MEM[1938] + MEM[9311];
assign MEM[14118] = MEM[1942] + MEM[3221];
assign MEM[14119] = MEM[1951] + MEM[4438];
assign MEM[14120] = MEM[1954] + MEM[2783];
assign MEM[14121] = MEM[1956] + MEM[9061];
assign MEM[14122] = MEM[1959] + MEM[2530];
assign MEM[14123] = MEM[1962] + MEM[5947];
assign MEM[14124] = MEM[1966] + MEM[3450];
assign MEM[14125] = MEM[1967] + MEM[2100];
assign MEM[14126] = MEM[1978] + MEM[6722];
assign MEM[14127] = MEM[1980] + MEM[4183];
assign MEM[14128] = MEM[1981] + MEM[463];
assign MEM[14129] = MEM[1988] + MEM[5525];
assign MEM[14130] = MEM[1996] + MEM[2151];
assign MEM[14131] = MEM[2015] + MEM[13503];
assign MEM[14132] = MEM[2021] + MEM[6899];
assign MEM[14133] = MEM[2022] + MEM[1255];
assign MEM[14134] = MEM[2022] + MEM[8190];
assign MEM[14135] = MEM[2031] + MEM[2679];
assign MEM[14136] = MEM[2037] + MEM[3053];
assign MEM[14137] = MEM[2039] + MEM[9278];
assign MEM[14138] = MEM[2043] + MEM[7025];
assign MEM[14139] = MEM[2050] + MEM[3034];
assign MEM[14140] = MEM[2055] + MEM[3263];
assign MEM[14141] = MEM[2058] + MEM[5332];
assign MEM[14142] = MEM[2069] + MEM[2581];
assign MEM[14143] = MEM[2087] + MEM[3941];
assign MEM[14144] = MEM[2090] + MEM[7926];
assign MEM[14145] = MEM[2091] + MEM[2309];
assign MEM[14146] = MEM[2099] + MEM[8863];
assign MEM[14147] = MEM[2102] + MEM[6571];
assign MEM[14148] = MEM[2108] + MEM[3682];
assign MEM[14149] = MEM[2114] + MEM[9745];
assign MEM[14150] = MEM[2125] + MEM[5407];
assign MEM[14151] = MEM[2143] + MEM[3787];
assign MEM[14152] = MEM[2166] + MEM[4974];
assign MEM[14153] = MEM[2170] + MEM[4911];
assign MEM[14154] = MEM[2178] + MEM[5190];
assign MEM[14155] = MEM[2186] + MEM[4599];
assign MEM[14156] = MEM[2195] + MEM[2294];
assign MEM[14157] = MEM[2197] + MEM[2834];
assign MEM[14158] = MEM[2202] + MEM[2436];
assign MEM[14159] = MEM[2203] + MEM[6893];
assign MEM[14160] = MEM[2212] + MEM[8244];
assign MEM[14161] = MEM[2218] + MEM[5101];
assign MEM[14162] = MEM[2220] + MEM[6134];
assign MEM[14163] = MEM[2226] + MEM[3901];
assign MEM[14164] = MEM[2231] + MEM[4463];
assign MEM[14165] = MEM[2254] + MEM[1108];
assign MEM[14166] = MEM[2278] + MEM[4927];
assign MEM[14167] = MEM[2287] + MEM[4934];
assign MEM[14168] = MEM[2291] + MEM[6317];
assign MEM[14169] = MEM[2295] + MEM[5363];
assign MEM[14170] = MEM[2301] + MEM[1898];
assign MEM[14171] = MEM[2308] + MEM[2629];
assign MEM[14172] = MEM[2315] + MEM[7204];
assign MEM[14173] = MEM[2331] + MEM[8706];
assign MEM[14174] = MEM[2333] + MEM[9057];
assign MEM[14175] = MEM[2334] + MEM[2674];
assign MEM[14176] = MEM[2335] + MEM[3842];
assign MEM[14177] = MEM[2338] + MEM[2673];
assign MEM[14178] = MEM[2339] + MEM[7467];
assign MEM[14179] = MEM[2348] + MEM[3284];
assign MEM[14180] = MEM[2349] + MEM[7385];
assign MEM[14181] = MEM[2351] + MEM[7322];
assign MEM[14182] = MEM[2356] + MEM[8557];
assign MEM[14183] = MEM[2359] + MEM[5706];
assign MEM[14184] = MEM[2367] + MEM[11212];
assign MEM[14185] = MEM[2374] + MEM[8595];
assign MEM[14186] = MEM[2379] + MEM[7560];
assign MEM[14187] = MEM[2389] + MEM[7042];
assign MEM[14188] = MEM[2413] + MEM[5911];
assign MEM[14189] = MEM[2415] + MEM[5166];
assign MEM[14190] = MEM[2421] + MEM[2854];
assign MEM[14191] = MEM[2422] + MEM[5422];
assign MEM[14192] = MEM[2452] + MEM[3573];
assign MEM[14193] = MEM[2455] + MEM[2893];
assign MEM[14194] = MEM[2482] + MEM[5158];
assign MEM[14195] = MEM[2485] + MEM[7271];
assign MEM[14196] = MEM[2487] + MEM[2749];
assign MEM[14197] = MEM[2492] + MEM[10154];
assign MEM[14198] = MEM[2503] + MEM[2718];
assign MEM[14199] = MEM[2514] + MEM[2885];
assign MEM[14200] = MEM[2517] + MEM[7354];
assign MEM[14201] = MEM[2523] + MEM[7712];
assign MEM[14202] = MEM[2525] + MEM[2951];
assign MEM[14203] = MEM[2526] + MEM[4157];
assign MEM[14204] = MEM[2527] + MEM[3090];
assign MEM[14205] = MEM[2539] + MEM[4803];
assign MEM[14206] = MEM[2556] + MEM[3117];
assign MEM[14207] = MEM[2567] + MEM[7516];
assign MEM[14208] = MEM[2570] + MEM[5870];
assign MEM[14209] = MEM[2578] + MEM[4150];
assign MEM[14210] = MEM[2582] + MEM[7702];
assign MEM[14211] = MEM[2583] + MEM[5195];
assign MEM[14212] = MEM[2588] + MEM[6548];
assign MEM[14213] = MEM[2589] + MEM[10896];
assign MEM[14214] = MEM[2590] + MEM[6276];
assign MEM[14215] = MEM[2591] + MEM[7908];
assign MEM[14216] = MEM[2598] + MEM[4269];
assign MEM[14217] = MEM[2603] + MEM[7503];
assign MEM[14218] = MEM[2604] + MEM[8420];
assign MEM[14219] = MEM[2610] + MEM[7127];
assign MEM[14220] = MEM[2611] + MEM[8386];
assign MEM[14221] = MEM[2614] + MEM[5133];
assign MEM[14222] = MEM[2622] + MEM[6370];
assign MEM[14223] = MEM[2644] + MEM[7069];
assign MEM[14224] = MEM[2647] + MEM[4134];
assign MEM[14225] = MEM[2651] + MEM[8296];
assign MEM[14226] = MEM[2655] + MEM[3859];
assign MEM[14227] = MEM[2658] + MEM[3781];
assign MEM[14228] = MEM[2660] + MEM[7870];
assign MEM[14229] = MEM[2662] + MEM[8465];
assign MEM[14230] = MEM[2668] + MEM[4642];
assign MEM[14231] = MEM[2671] + MEM[3725];
assign MEM[14232] = MEM[2678] + MEM[2823];
assign MEM[14233] = MEM[2692] + MEM[3082];
assign MEM[14234] = MEM[2693] + MEM[6341];
assign MEM[14235] = MEM[2694] + MEM[5110];
assign MEM[14236] = MEM[2699] + MEM[3124];
assign MEM[14237] = MEM[2703] + MEM[7986];
assign MEM[14238] = MEM[2722] + MEM[7985];
assign MEM[14239] = MEM[2726] + MEM[8556];
assign MEM[14240] = MEM[2727] + MEM[6182];
assign MEM[14241] = MEM[2730] + MEM[4627];
assign MEM[14242] = MEM[2743] + MEM[6124];
assign MEM[14243] = MEM[2747] + MEM[8428];
assign MEM[14244] = MEM[2754] + MEM[7793];
assign MEM[14245] = MEM[2757] + MEM[3270];
assign MEM[14246] = MEM[2762] + MEM[4531];
assign MEM[14247] = MEM[2765] + MEM[5866];
assign MEM[14248] = MEM[2773] + MEM[7609];
assign MEM[14249] = MEM[2774] + MEM[3126];
assign MEM[14250] = MEM[2780] + MEM[4621];
assign MEM[14251] = MEM[2781] + MEM[4454];
assign MEM[14252] = MEM[2791] + MEM[3388];
assign MEM[14253] = MEM[2797] + MEM[9088];
assign MEM[14254] = MEM[2802] + MEM[5758];
assign MEM[14255] = MEM[2810] + MEM[4268];
assign MEM[14256] = MEM[2826] + MEM[8204];
assign MEM[14257] = MEM[2843] + MEM[10758];
assign MEM[14258] = MEM[2850] + MEM[5695];
assign MEM[14259] = MEM[2855] + MEM[8490];
assign MEM[14260] = MEM[2867] + MEM[3415];
assign MEM[14261] = MEM[2868] + MEM[9617];
assign MEM[14262] = MEM[2874] + MEM[8849];
assign MEM[14263] = MEM[2876] + MEM[9355];
assign MEM[14264] = MEM[2877] + MEM[7429];
assign MEM[14265] = MEM[2878] + MEM[5891];
assign MEM[14266] = MEM[2878] + MEM[11566];
assign MEM[14267] = MEM[2890] + MEM[8914];
assign MEM[14268] = MEM[2898] + MEM[3007];
assign MEM[14269] = MEM[2898] + MEM[10787];
assign MEM[14270] = MEM[2900] + MEM[7875];
assign MEM[14271] = MEM[2932] + MEM[6345];
assign MEM[14272] = MEM[2938] + MEM[4230];
assign MEM[14273] = MEM[2948] + MEM[8717];
assign MEM[14274] = MEM[2962] + MEM[5338];
assign MEM[14275] = MEM[2966] + MEM[7477];
assign MEM[14276] = MEM[2970] + MEM[5670];
assign MEM[14277] = MEM[2975] + MEM[7549];
assign MEM[14278] = MEM[2979] + MEM[7540];
assign MEM[14279] = MEM[2980] + MEM[3076];
assign MEM[14280] = MEM[2988] + MEM[3299];
assign MEM[14281] = MEM[2990] + MEM[4851];
assign MEM[14282] = MEM[2997] + MEM[8293];
assign MEM[14283] = MEM[3011] + MEM[9721];
assign MEM[14284] = MEM[3018] + MEM[8509];
assign MEM[14285] = MEM[3021] + MEM[3797];
assign MEM[14286] = MEM[3027] + MEM[8314];
assign MEM[14287] = MEM[3028] + MEM[4998];
assign MEM[14288] = MEM[3036] + MEM[5540];
assign MEM[14289] = MEM[3061] + MEM[6937];
assign MEM[14290] = MEM[3066] + MEM[7787];
assign MEM[14291] = MEM[3086] + MEM[3851];
assign MEM[14292] = MEM[3093] + MEM[8186];
assign MEM[14293] = MEM[3106] + MEM[3235];
assign MEM[14294] = MEM[3107] + MEM[9965];
assign MEM[14295] = MEM[3116] + MEM[4019];
assign MEM[14296] = MEM[3122] + MEM[7964];
assign MEM[14297] = MEM[3123] + MEM[3618];
assign MEM[14298] = MEM[3134] + MEM[3620];
assign MEM[14299] = MEM[3135] + MEM[5125];
assign MEM[14300] = MEM[3143] + MEM[6101];
assign MEM[14301] = MEM[3149] + MEM[8986];
assign MEM[14302] = MEM[3158] + MEM[5312];
assign MEM[14303] = MEM[3164] + MEM[4590];
assign MEM[14304] = MEM[3171] + MEM[4046];
assign MEM[14305] = MEM[3175] + MEM[7550];
assign MEM[14306] = MEM[3179] + MEM[3899];
assign MEM[14307] = MEM[3180] + MEM[5150];
assign MEM[14308] = MEM[3183] + MEM[8323];
assign MEM[14309] = MEM[3187] + MEM[7441];
assign MEM[14310] = MEM[3215] + MEM[5313];
assign MEM[14311] = MEM[3218] + MEM[4852];
assign MEM[14312] = MEM[3223] + MEM[8384];
assign MEM[14313] = MEM[3239] + MEM[9048];
assign MEM[14314] = MEM[3244] + MEM[3786];
assign MEM[14315] = MEM[3252] + MEM[10367];
assign MEM[14316] = MEM[3261] + MEM[9736];
assign MEM[14317] = MEM[3266] + MEM[9390];
assign MEM[14318] = MEM[3267] + MEM[7679];
assign MEM[14319] = MEM[3268] + MEM[3827];
assign MEM[14320] = MEM[3278] + MEM[7808];
assign MEM[14321] = MEM[3298] + MEM[4382];
assign MEM[14322] = MEM[3301] + MEM[6656];
assign MEM[14323] = MEM[3303] + MEM[6505];
assign MEM[14324] = MEM[3307] + MEM[4427];
assign MEM[14325] = MEM[3341] + MEM[4236];
assign MEM[14326] = MEM[3343] + MEM[7698];
assign MEM[14327] = MEM[3372] + MEM[7173];
assign MEM[14328] = MEM[3390] + MEM[4242];
assign MEM[14329] = MEM[3395] + MEM[8946];
assign MEM[14330] = MEM[3396] + MEM[3564];
assign MEM[14331] = MEM[3406] + MEM[9154];
assign MEM[14332] = MEM[3414] + MEM[3500];
assign MEM[14333] = MEM[3426] + MEM[7121];
assign MEM[14334] = MEM[3427] + MEM[6702];
assign MEM[14335] = MEM[3431] + MEM[4290];
assign MEM[14336] = MEM[3435] + MEM[7297];
assign MEM[14337] = MEM[3438] + MEM[8527];
assign MEM[14338] = MEM[3446] + MEM[8232];
assign MEM[14339] = MEM[3451] + MEM[7431];
assign MEM[14340] = MEM[3459] + MEM[4202];
assign MEM[14341] = MEM[3470] + MEM[8074];
assign MEM[14342] = MEM[3492] + MEM[5427];
assign MEM[14343] = MEM[3498] + MEM[8457];
assign MEM[14344] = MEM[3510] + MEM[4636];
assign MEM[14345] = MEM[3518] + MEM[6339];
assign MEM[14346] = MEM[3524] + MEM[4462];
assign MEM[14347] = MEM[3533] + MEM[7372];
assign MEM[14348] = MEM[3535] + MEM[6606];
assign MEM[14349] = MEM[3540] + MEM[5403];
assign MEM[14350] = MEM[3541] + MEM[5395];
assign MEM[14351] = MEM[3566] + MEM[4603];
assign MEM[14352] = MEM[3578] + MEM[7236];
assign MEM[14353] = MEM[3580] + MEM[7561];
assign MEM[14354] = MEM[3581] + MEM[10926];
assign MEM[14355] = MEM[3589] + MEM[5014];
assign MEM[14356] = MEM[3597] + MEM[8448];
assign MEM[14357] = MEM[3598] + MEM[7049];
assign MEM[14358] = MEM[3606] + MEM[8864];
assign MEM[14359] = MEM[3612] + MEM[7551];
assign MEM[14360] = MEM[3634] + MEM[4418];
assign MEM[14361] = MEM[3642] + MEM[8751];
assign MEM[14362] = MEM[3643] + MEM[3995];
assign MEM[14363] = MEM[3647] + MEM[8501];
assign MEM[14364] = MEM[3654] + MEM[8959];
assign MEM[14365] = MEM[3677] + MEM[4935];
assign MEM[14366] = MEM[3685] + MEM[5917];
assign MEM[14367] = MEM[3692] + MEM[5467];
assign MEM[14368] = MEM[3703] + MEM[8086];
assign MEM[14369] = MEM[3710] + MEM[7701];
assign MEM[14370] = MEM[3711] + MEM[8811];
assign MEM[14371] = MEM[3715] + MEM[10906];
assign MEM[14372] = MEM[3717] + MEM[8671];
assign MEM[14373] = MEM[3722] + MEM[4044];
assign MEM[14374] = MEM[3723] + MEM[6564];
assign MEM[14375] = MEM[3734] + MEM[7562];
assign MEM[14376] = MEM[3751] + MEM[3571];
assign MEM[14377] = MEM[3757] + MEM[9302];
assign MEM[14378] = MEM[3766] + MEM[11054];
assign MEM[14379] = MEM[3767] + MEM[5215];
assign MEM[14380] = MEM[3771] + MEM[8409];
assign MEM[14381] = MEM[3782] + MEM[5068];
assign MEM[14382] = MEM[3783] + MEM[8529];
assign MEM[14383] = MEM[3794] + MEM[5687];
assign MEM[14384] = MEM[3796] + MEM[8298];
assign MEM[14385] = MEM[3798] + MEM[6031];
assign MEM[14386] = MEM[3802] + MEM[6148];
assign MEM[14387] = MEM[3803] + MEM[5350];
assign MEM[14388] = MEM[3830] + MEM[7349];
assign MEM[14389] = MEM[3850] + MEM[9463];
assign MEM[14390] = MEM[3868] + MEM[6610];
assign MEM[14391] = MEM[3869] + MEM[5805];
assign MEM[14392] = MEM[3871] + MEM[4538];
assign MEM[14393] = MEM[3890] + MEM[7480];
assign MEM[14394] = MEM[3900] + MEM[9942];
assign MEM[14395] = MEM[3908] + MEM[7711];
assign MEM[14396] = MEM[3909] + MEM[8851];
assign MEM[14397] = MEM[3914] + MEM[5254];
assign MEM[14398] = MEM[3916] + MEM[4381];
assign MEM[14399] = MEM[3917] + MEM[6433];
assign MEM[14400] = MEM[3931] + MEM[7911];
assign MEM[14401] = MEM[3939] + MEM[8568];
assign MEM[14402] = MEM[3946] + MEM[7660];
assign MEM[14403] = MEM[3947] + MEM[6102];
assign MEM[14404] = MEM[3951] + MEM[8330];
assign MEM[14405] = MEM[3970] + MEM[4970];
assign MEM[14406] = MEM[3974] + MEM[7547];
assign MEM[14407] = MEM[3975] + MEM[5763];
assign MEM[14408] = MEM[3997] + MEM[8304];
assign MEM[14409] = MEM[4007] + MEM[5666];
assign MEM[14410] = MEM[4010] + MEM[9005];
assign MEM[14411] = MEM[4012] + MEM[10073];
assign MEM[14412] = MEM[4039] + MEM[4855];
assign MEM[14413] = MEM[4045] + MEM[6478];
assign MEM[14414] = MEM[4055] + MEM[7644];
assign MEM[14415] = MEM[4063] + MEM[7771];
assign MEM[14416] = MEM[4070] + MEM[6255];
assign MEM[14417] = MEM[4085] + MEM[8138];
assign MEM[14418] = MEM[4107] + MEM[8470];
assign MEM[14419] = MEM[4109] + MEM[6188];
assign MEM[14420] = MEM[4119] + MEM[5692];
assign MEM[14421] = MEM[4133] + MEM[5198];
assign MEM[14422] = MEM[4178] + MEM[9291];
assign MEM[14423] = MEM[4179] + MEM[10940];
assign MEM[14424] = MEM[4181] + MEM[7035];
assign MEM[14425] = MEM[4182] + MEM[7491];
assign MEM[14426] = MEM[4183] + MEM[8940];
assign MEM[14427] = MEM[4195] + MEM[5750];
assign MEM[14428] = MEM[4203] + MEM[9760];
assign MEM[14429] = MEM[4212] + MEM[6213];
assign MEM[14430] = MEM[4227] + MEM[4534];
assign MEM[14431] = MEM[4234] + MEM[6674];
assign MEM[14432] = MEM[4244] + MEM[8432];
assign MEM[14433] = MEM[4270] + MEM[4539];
assign MEM[14434] = MEM[4276] + MEM[4429];
assign MEM[14435] = MEM[4279] + MEM[8160];
assign MEM[14436] = MEM[4284] + MEM[10752];
assign MEM[14437] = MEM[4299] + MEM[6011];
assign MEM[14438] = MEM[4302] + MEM[4892];
assign MEM[14439] = MEM[4310] + MEM[6555];
assign MEM[14440] = MEM[4311] + MEM[6871];
assign MEM[14441] = MEM[4323] + MEM[5402];
assign MEM[14442] = MEM[4332] + MEM[8396];
assign MEM[14443] = MEM[4334] + MEM[4989];
assign MEM[14444] = MEM[4354] + MEM[7871];
assign MEM[14445] = MEM[4364] + MEM[7410];
assign MEM[14446] = MEM[4371] + MEM[5821];
assign MEM[14447] = MEM[4372] + MEM[6330];
assign MEM[14448] = MEM[4380] + MEM[5988];
assign MEM[14449] = MEM[4386] + MEM[8510];
assign MEM[14450] = MEM[4396] + MEM[8605];
assign MEM[14451] = MEM[4403] + MEM[2972];
assign MEM[14452] = MEM[4404] + MEM[7643];
assign MEM[14453] = MEM[4421] + MEM[5455];
assign MEM[14454] = MEM[4422] + MEM[9515];
assign MEM[14455] = MEM[4428] + MEM[9966];
assign MEM[14456] = MEM[4434] + MEM[8239];
assign MEM[14457] = MEM[4438] + MEM[9699];
assign MEM[14458] = MEM[4445] + MEM[5181];
assign MEM[14459] = MEM[4458] + MEM[8461];
assign MEM[14460] = MEM[4459] + MEM[6294];
assign MEM[14461] = MEM[4467] + MEM[5197];
assign MEM[14462] = MEM[4468] + MEM[2403];
assign MEM[14463] = MEM[4471] + MEM[8176];
assign MEM[14464] = MEM[4475] + MEM[10021];
assign MEM[14465] = MEM[4476] + MEM[7118];
assign MEM[14466] = MEM[4479] + MEM[6157];
assign MEM[14467] = MEM[4486] + MEM[7859];
assign MEM[14468] = MEM[4491] + MEM[6778];
assign MEM[14469] = MEM[4492] + MEM[5767];
assign MEM[14470] = MEM[4494] + MEM[10703];
assign MEM[14471] = MEM[4500] + MEM[6150];
assign MEM[14472] = MEM[4514] + MEM[9979];
assign MEM[14473] = MEM[4518] + MEM[5309];
assign MEM[14474] = MEM[4523] + MEM[8804];
assign MEM[14475] = MEM[4526] + MEM[6245];
assign MEM[14476] = MEM[4541] + MEM[7119];
assign MEM[14477] = MEM[4547] + MEM[6697];
assign MEM[14478] = MEM[4551] + MEM[9960];
assign MEM[14479] = MEM[4572] + MEM[10040];
assign MEM[14480] = MEM[4620] + MEM[7854];
assign MEM[14481] = MEM[4622] + MEM[7910];
assign MEM[14482] = MEM[4628] + MEM[7536];
assign MEM[14483] = MEM[4634] + MEM[8277];
assign MEM[14484] = MEM[4637] + MEM[9913];
assign MEM[14485] = MEM[4643] + MEM[10037];
assign MEM[14486] = MEM[4651] + MEM[4767];
assign MEM[14487] = MEM[4662] + MEM[5639];
assign MEM[14488] = MEM[4663] + MEM[9410];
assign MEM[14489] = MEM[4678] + MEM[9293];
assign MEM[14490] = MEM[4684] + MEM[6464];
assign MEM[14491] = MEM[4685] + MEM[10754];
assign MEM[14492] = MEM[4691] + MEM[9527];
assign MEM[14493] = MEM[4694] + MEM[9203];
assign MEM[14494] = MEM[4702] + MEM[8361];
assign MEM[14495] = MEM[4719] + MEM[8885];
assign MEM[14496] = MEM[4749] + MEM[7707];
assign MEM[14497] = MEM[4755] + MEM[6506];
assign MEM[14498] = MEM[4756] + MEM[8078];
assign MEM[14499] = MEM[4757] + MEM[4780];
assign MEM[14500] = MEM[4758] + MEM[9855];
assign MEM[14501] = MEM[4759] + MEM[10772];
assign MEM[14502] = MEM[4771] + MEM[3805];
assign MEM[14503] = MEM[4772] + MEM[7508];
assign MEM[14504] = MEM[4774] + MEM[10931];
assign MEM[14505] = MEM[4789] + MEM[6140];
assign MEM[14506] = MEM[4810] + MEM[4887];
assign MEM[14507] = MEM[4814] + MEM[8071];
assign MEM[14508] = MEM[4823] + MEM[10308];
assign MEM[14509] = MEM[4836] + MEM[7455];
assign MEM[14510] = MEM[4854] + MEM[9893];
assign MEM[14511] = MEM[4859] + MEM[8162];
assign MEM[14512] = MEM[4863] + MEM[5860];
assign MEM[14513] = MEM[4868] + MEM[6523];
assign MEM[14514] = MEM[4882] + MEM[8214];
assign MEM[14515] = MEM[4893] + MEM[8693];
assign MEM[14516] = MEM[4898] + MEM[11087];
assign MEM[14517] = MEM[4899] + MEM[8581];
assign MEM[14518] = MEM[4949] + MEM[7662];
assign MEM[14519] = MEM[4955] + MEM[8526];
assign MEM[14520] = MEM[4956] + MEM[6799];
assign MEM[14521] = MEM[4965] + MEM[7913];
assign MEM[14522] = MEM[4971] + MEM[7747];
assign MEM[14523] = MEM[4974] + MEM[8262];
assign MEM[14524] = MEM[4978] + MEM[5562];
assign MEM[14525] = MEM[4986] + MEM[6434];
assign MEM[14526] = MEM[4990] + MEM[7395];
assign MEM[14527] = MEM[5005] + MEM[7675];
assign MEM[14528] = MEM[5011] + MEM[9957];
assign MEM[14529] = MEM[5019] + MEM[5659];
assign MEM[14530] = MEM[5023] + MEM[5443];
assign MEM[14531] = MEM[5042] + MEM[9120];
assign MEM[14532] = MEM[5050] + MEM[7561];
assign MEM[14533] = MEM[5061] + MEM[8399];
assign MEM[14534] = MEM[5086] + MEM[8727];
assign MEM[14535] = MEM[5106] + MEM[6085];
assign MEM[14536] = MEM[5118] + MEM[7745];
assign MEM[14537] = MEM[5132] + MEM[10304];
assign MEM[14538] = MEM[5139] + MEM[8476];
assign MEM[14539] = MEM[5149] + MEM[7989];
assign MEM[14540] = MEM[5157] + MEM[6187];
assign MEM[14541] = MEM[5172] + MEM[6438];
assign MEM[14542] = MEM[5189] + MEM[7152];
assign MEM[14543] = MEM[5205] + MEM[3403];
assign MEM[14544] = MEM[5218] + MEM[7813];
assign MEM[14545] = MEM[5219] + MEM[7442];
assign MEM[14546] = MEM[5221] + MEM[8192];
assign MEM[14547] = MEM[5230] + MEM[8254];
assign MEM[14548] = MEM[5236] + MEM[8141];
assign MEM[14549] = MEM[5286] + MEM[8560];
assign MEM[14550] = MEM[5326] + MEM[7478];
assign MEM[14551] = MEM[5343] + MEM[8917];
assign MEM[14552] = MEM[5346] + MEM[3879];
assign MEM[14553] = MEM[5348] + MEM[9220];
assign MEM[14554] = MEM[5349] + MEM[7326];
assign MEM[14555] = MEM[5357] + MEM[7369];
assign MEM[14556] = MEM[5375] + MEM[1670];
assign MEM[14557] = MEM[5434] + MEM[6375];
assign MEM[14558] = MEM[5447] + MEM[8523];
assign MEM[14559] = MEM[5450] + MEM[10053];
assign MEM[14560] = MEM[5468] + MEM[8801];
assign MEM[14561] = MEM[5477] + MEM[9083];
assign MEM[14562] = MEM[5478] + MEM[7881];
assign MEM[14563] = MEM[5479] + MEM[6334];
assign MEM[14564] = MEM[5507] + MEM[8098];
assign MEM[14565] = MEM[5542] + MEM[6662];
assign MEM[14566] = MEM[5543] + MEM[7352];
assign MEM[14567] = MEM[5549] + MEM[7785];
assign MEM[14568] = MEM[5582] + MEM[7725];
assign MEM[14569] = MEM[5605] + MEM[9379];
assign MEM[14570] = MEM[5645] + MEM[10460];
assign MEM[14571] = MEM[5647] + MEM[10197];
assign MEM[14572] = MEM[5651] + MEM[8131];
assign MEM[14573] = MEM[5653] + MEM[6737];
assign MEM[14574] = MEM[5658] + MEM[8064];
assign MEM[14575] = MEM[5675] + MEM[9450];
assign MEM[14576] = MEM[5676] + MEM[7367];
assign MEM[14577] = MEM[5677] + MEM[7915];
assign MEM[14578] = MEM[5683] + MEM[7933];
assign MEM[14579] = MEM[5693] + MEM[8780];
assign MEM[14580] = MEM[5698] + MEM[8030];
assign MEM[14581] = MEM[5699] + MEM[10882];
assign MEM[14582] = MEM[5709] + MEM[8668];
assign MEM[14583] = MEM[5723] + MEM[5885];
assign MEM[14584] = MEM[5737] + MEM[8473];
assign MEM[14585] = MEM[5739] + MEM[8164];
assign MEM[14586] = MEM[5740] + MEM[6215];
assign MEM[14587] = MEM[5743] + MEM[8415];
assign MEM[14588] = MEM[5775] + MEM[5708];
assign MEM[14589] = MEM[5789] + MEM[8187];
assign MEM[14590] = MEM[5795] + MEM[8210];
assign MEM[14591] = MEM[5806] + MEM[7535];
assign MEM[14592] = MEM[5831] + MEM[6618];
assign MEM[14593] = MEM[5837] + MEM[10688];
assign MEM[14594] = MEM[5862] + MEM[6253];
assign MEM[14595] = MEM[5876] + MEM[8143];
assign MEM[14596] = MEM[5884] + MEM[8280];
assign MEM[14597] = MEM[5886] + MEM[2274];
assign MEM[14598] = MEM[5894] + MEM[3466];
assign MEM[14599] = MEM[5896] + MEM[8216];
assign MEM[14600] = MEM[5897] + MEM[9848];
assign MEM[14601] = MEM[5954] + MEM[9039];
assign MEM[14602] = MEM[5965] + MEM[6516];
assign MEM[14603] = MEM[5995] + MEM[6605];
assign MEM[14604] = MEM[6006] + MEM[8130];
assign MEM[14605] = MEM[6007] + MEM[7499];
assign MEM[14606] = MEM[6013] + MEM[8261];
assign MEM[14607] = MEM[6030] + MEM[8732];
assign MEM[14608] = MEM[6079] + MEM[7389];
assign MEM[14609] = MEM[6109] + MEM[9858];
assign MEM[14610] = MEM[6110] + MEM[6836];
assign MEM[14611] = MEM[6126] + MEM[4580];
assign MEM[14612] = MEM[6139] + MEM[10042];
assign MEM[14613] = MEM[6147] + MEM[8737];
assign MEM[14614] = MEM[6181] + MEM[6322];
assign MEM[14615] = MEM[6219] + MEM[8482];
assign MEM[14616] = MEM[6222] + MEM[6254];
assign MEM[14617] = MEM[6223] + MEM[9959];
assign MEM[14618] = MEM[6227] + MEM[8749];
assign MEM[14619] = MEM[6228] + MEM[7539];
assign MEM[14620] = MEM[6245] + MEM[9289];
assign MEM[14621] = MEM[6247] + MEM[8785];
assign MEM[14622] = MEM[6255] + MEM[10928];
assign MEM[14623] = MEM[6284] + MEM[8349];
assign MEM[14624] = MEM[6290] + MEM[10898];
assign MEM[14625] = MEM[6302] + MEM[7548];
assign MEM[14626] = MEM[6331] + MEM[9126];
assign MEM[14627] = MEM[6333] + MEM[939];
assign MEM[14628] = MEM[6338] + MEM[10853];
assign MEM[14629] = MEM[6340] + MEM[8335];
assign MEM[14630] = MEM[6344] + MEM[8365];
assign MEM[14631] = MEM[6359] + MEM[7756];
assign MEM[14632] = MEM[6366] + MEM[9183];
assign MEM[14633] = MEM[6377] + MEM[8844];
assign MEM[14634] = MEM[6402] + MEM[6613];
assign MEM[14635] = MEM[6405] + MEM[7869];
assign MEM[14636] = MEM[6410] + MEM[8255];
assign MEM[14637] = MEM[6420] + MEM[9811];
assign MEM[14638] = MEM[6425] + MEM[8484];
assign MEM[14639] = MEM[6428] + MEM[6997];
assign MEM[14640] = MEM[6442] + MEM[8621];
assign MEM[14641] = MEM[6472] + MEM[7975];
assign MEM[14642] = MEM[6485] + MEM[8155];
assign MEM[14643] = MEM[6490] + MEM[8610];
assign MEM[14644] = MEM[6496] + MEM[9219];
assign MEM[14645] = MEM[6497] + MEM[8497];
assign MEM[14646] = MEM[6501] + MEM[8888];
assign MEM[14647] = MEM[6517] + MEM[10328];
assign MEM[14648] = MEM[6546] + MEM[7733];
assign MEM[14649] = MEM[6557] + MEM[9119];
assign MEM[14650] = MEM[6562] + MEM[7339];
assign MEM[14651] = MEM[6566] + MEM[7468];
assign MEM[14652] = MEM[6577] + MEM[7000];
assign MEM[14653] = MEM[6581] + MEM[7281];
assign MEM[14654] = MEM[6583] + MEM[7315];
assign MEM[14655] = MEM[6585] + MEM[8100];
assign MEM[14656] = MEM[6593] + MEM[8072];
assign MEM[14657] = MEM[6598] + MEM[8992];
assign MEM[14658] = MEM[6612] + MEM[7970];
assign MEM[14659] = MEM[6631] + MEM[378];
assign MEM[14660] = MEM[6634] + MEM[10916];
assign MEM[14661] = MEM[6635] + MEM[8591];
assign MEM[14662] = MEM[6648] + MEM[9391];
assign MEM[14663] = MEM[6650] + MEM[9143];
assign MEM[14664] = MEM[6657] + MEM[7743];
assign MEM[14665] = MEM[6668] + MEM[6672];
assign MEM[14666] = MEM[6695] + MEM[7694];
assign MEM[14667] = MEM[6696] + MEM[7384];
assign MEM[14668] = MEM[6704] + MEM[11693];
assign MEM[14669] = MEM[6707] + MEM[7765];
assign MEM[14670] = MEM[6716] + MEM[7318];
assign MEM[14671] = MEM[6724] + MEM[10189];
assign MEM[14672] = MEM[6736] + MEM[7718];
assign MEM[14673] = MEM[6750] + MEM[10984];
assign MEM[14674] = MEM[6796] + MEM[7095];
assign MEM[14675] = MEM[6809] + MEM[9826];
assign MEM[14676] = MEM[6815] + MEM[8652];
assign MEM[14677] = MEM[6817] + MEM[7099];
assign MEM[14678] = MEM[6848] + MEM[8017];
assign MEM[14679] = MEM[6866] + MEM[6973];
assign MEM[14680] = MEM[6874] + MEM[7629];
assign MEM[14681] = MEM[6885] + MEM[8307];
assign MEM[14682] = MEM[6889] + MEM[8687];
assign MEM[14683] = MEM[6895] + MEM[9810];
assign MEM[14684] = MEM[6896] + MEM[8782];
assign MEM[14685] = MEM[6910] + MEM[7541];
assign MEM[14686] = MEM[6911] + MEM[9253];
assign MEM[14687] = MEM[6912] + MEM[8905];
assign MEM[14688] = MEM[6929] + MEM[7993];
assign MEM[14689] = MEM[6931] + MEM[9446];
assign MEM[14690] = MEM[6932] + MEM[8502];
assign MEM[14691] = MEM[6933] + MEM[10999];
assign MEM[14692] = MEM[6941] + MEM[8205];
assign MEM[14693] = MEM[6944] + MEM[8661];
assign MEM[14694] = MEM[6950] + MEM[7802];
assign MEM[14695] = MEM[6952] + MEM[8434];
assign MEM[14696] = MEM[6953] + MEM[9485];
assign MEM[14697] = MEM[6955] + MEM[8900];
assign MEM[14698] = MEM[6961] + MEM[11171];
assign MEM[14699] = MEM[6963] + MEM[8909];
assign MEM[14700] = MEM[6971] + MEM[8309];
assign MEM[14701] = MEM[6981] + MEM[8228];
assign MEM[14702] = MEM[6986] + MEM[7419];
assign MEM[14703] = MEM[6987] + MEM[8006];
assign MEM[14704] = MEM[6988] + MEM[9087];
assign MEM[14705] = MEM[6993] + MEM[6364];
assign MEM[14706] = MEM[7005] + MEM[8360];
assign MEM[14707] = MEM[7016] + MEM[9230];
assign MEM[14708] = MEM[7022] + MEM[9921];
assign MEM[14709] = MEM[7034] + MEM[7735];
assign MEM[14710] = MEM[7056] + MEM[7172];
assign MEM[14711] = MEM[7065] + MEM[8161];
assign MEM[14712] = MEM[7089] + MEM[9272];
assign MEM[14713] = MEM[7091] + MEM[10909];
assign MEM[14714] = MEM[7094] + MEM[8602];
assign MEM[14715] = MEM[7097] + MEM[2534];
assign MEM[14716] = MEM[7109] + MEM[9242];
assign MEM[14717] = MEM[7110] + MEM[9718];
assign MEM[14718] = MEM[7111] + MEM[8907];
assign MEM[14719] = MEM[7115] + MEM[7618];
assign MEM[14720] = MEM[7169] + MEM[7458];
assign MEM[14721] = MEM[7170] + MEM[7940];
assign MEM[14722] = MEM[7193] + MEM[8163];
assign MEM[14723] = MEM[7200] + MEM[9001];
assign MEM[14724] = MEM[7206] + MEM[7041];
assign MEM[14725] = MEM[7219] + MEM[9951];
assign MEM[14726] = MEM[7245] + MEM[7262];
assign MEM[14727] = MEM[7254] + MEM[10952];
assign MEM[14728] = MEM[7277] + MEM[7534];
assign MEM[14729] = MEM[7298] + MEM[7535];
assign MEM[14730] = MEM[7323] + MEM[7709];
assign MEM[14731] = MEM[7325] + MEM[8472];
assign MEM[14732] = MEM[7327] + MEM[9170];
assign MEM[14733] = MEM[7334] + MEM[8526];
assign MEM[14734] = MEM[7358] + MEM[10870];
assign MEM[14735] = MEM[7364] + MEM[8368];
assign MEM[14736] = MEM[7371] + MEM[8241];
assign MEM[14737] = MEM[7372] + MEM[8275];
assign MEM[14738] = MEM[7374] + MEM[8117];
assign MEM[14739] = MEM[7420] + MEM[8910];
assign MEM[14740] = MEM[7422] + MEM[8752];
assign MEM[14741] = MEM[7424] + MEM[8609];
assign MEM[14742] = MEM[7436] + MEM[4795];
assign MEM[14743] = MEM[7451] + MEM[7973];
assign MEM[14744] = MEM[7452] + MEM[8520];
assign MEM[14745] = MEM[7457] + MEM[7820];
assign MEM[14746] = MEM[7471] + MEM[8418];
assign MEM[14747] = MEM[7472] + MEM[8289];
assign MEM[14748] = MEM[7486] + MEM[10788];
assign MEM[14749] = MEM[7495] + MEM[9448];
assign MEM[14750] = MEM[7497] + MEM[8090];
assign MEM[14751] = MEM[7510] + MEM[8644];
assign MEM[14752] = MEM[7518] + MEM[8892];
assign MEM[14753] = MEM[7523] + MEM[8425];
assign MEM[14754] = MEM[7524] + MEM[3102];
assign MEM[14755] = MEM[7545] + MEM[10210];
assign MEM[14756] = MEM[7547] + MEM[8753];
assign MEM[14757] = MEM[7552] + MEM[7994];
assign MEM[14758] = MEM[7576] + MEM[8793];
assign MEM[14759] = MEM[7589] + MEM[8674];
assign MEM[14760] = MEM[7595] + MEM[8004];
assign MEM[14761] = MEM[7601] + MEM[7684];
assign MEM[14762] = MEM[7605] + MEM[8332];
assign MEM[14763] = MEM[7616] + MEM[8708];
assign MEM[14764] = MEM[7633] + MEM[9185];
assign MEM[14765] = MEM[7646] + MEM[8604];
assign MEM[14766] = MEM[7648] + MEM[9283];
assign MEM[14767] = MEM[7651] + MEM[11494];
assign MEM[14768] = MEM[7673] + MEM[8783];
assign MEM[14769] = MEM[7676] + MEM[8001];
assign MEM[14770] = MEM[7677] + MEM[582];
assign MEM[14771] = MEM[7690] + MEM[9539];
assign MEM[14772] = MEM[7702] + MEM[11234];
assign MEM[14773] = MEM[7704] + MEM[8059];
assign MEM[14774] = MEM[7723] + MEM[9031];
assign MEM[14775] = MEM[7724] + MEM[11241];
assign MEM[14776] = MEM[7727] + MEM[8250];
assign MEM[14777] = MEM[7731] + MEM[8957];
assign MEM[14778] = MEM[7739] + MEM[10929];
assign MEM[14779] = MEM[7746] + MEM[9103];
assign MEM[14780] = MEM[7761] + MEM[8125];
assign MEM[14781] = MEM[7770] + MEM[8555];
assign MEM[14782] = MEM[7789] + MEM[10153];
assign MEM[14783] = MEM[7791] + MEM[726];
assign MEM[14784] = MEM[7795] + MEM[11107];
assign MEM[14785] = MEM[7804] + MEM[8587];
assign MEM[14786] = MEM[7824] + MEM[8865];
assign MEM[14787] = MEM[7827] + MEM[1005];
assign MEM[14788] = MEM[7836] + MEM[9271];
assign MEM[14789] = MEM[7841] + MEM[9375];
assign MEM[14790] = MEM[7850] + MEM[6673];
assign MEM[14791] = MEM[7850] + MEM[10147];
assign MEM[14792] = MEM[7852] + MEM[8803];
assign MEM[14793] = MEM[7858] + MEM[8802];
assign MEM[14794] = MEM[7862] + MEM[2060];
assign MEM[14795] = MEM[7883] + MEM[7914];
assign MEM[14796] = MEM[7887] + MEM[9781];
assign MEM[14797] = MEM[7890] + MEM[8199];
assign MEM[14798] = MEM[7891] + MEM[9268];
assign MEM[14799] = MEM[7897] + MEM[8463];
assign MEM[14800] = MEM[7918] + MEM[8876];
assign MEM[14801] = MEM[7919] + MEM[8382];
assign MEM[14802] = MEM[7927] + MEM[9142];
assign MEM[14803] = MEM[7931] + MEM[8584];
assign MEM[14804] = MEM[7944] + MEM[8052];
assign MEM[14805] = MEM[7945] + MEM[8977];
assign MEM[14806] = MEM[7946] + MEM[8566];
assign MEM[14807] = MEM[7947] + MEM[6167];
assign MEM[14808] = MEM[7948] + MEM[8225];
assign MEM[14809] = MEM[7949] + MEM[8460];
assign MEM[14810] = MEM[7952] + MEM[9350];
assign MEM[14811] = MEM[7965] + MEM[9441];
assign MEM[14812] = MEM[8000] + MEM[10859];
assign MEM[14813] = MEM[8005] + MEM[10547];
assign MEM[14814] = MEM[8007] + MEM[2519];
assign MEM[14815] = MEM[8009] + MEM[9437];
assign MEM[14816] = MEM[8012] + MEM[6613];
assign MEM[14817] = MEM[8014] + MEM[8531];
assign MEM[14818] = MEM[8016] + MEM[8223];
assign MEM[14819] = MEM[8018] + MEM[8107];
assign MEM[14820] = MEM[8022] + MEM[9274];
assign MEM[14821] = MEM[8023] + MEM[9784];
assign MEM[14822] = MEM[8029] + MEM[8891];
assign MEM[14823] = MEM[8031] + MEM[8238];
assign MEM[14824] = MEM[8033] + MEM[8426];
assign MEM[14825] = MEM[8035] + MEM[8110];
assign MEM[14826] = MEM[8037] + MEM[9387];
assign MEM[14827] = MEM[8041] + MEM[9236];
assign MEM[14828] = MEM[8044] + MEM[7865];
assign MEM[14829] = MEM[8046] + MEM[7882];
assign MEM[14830] = MEM[8051] + MEM[5282];
assign MEM[14831] = MEM[8079] + MEM[11064];
assign MEM[14832] = MEM[8103] + MEM[8268];
assign MEM[14833] = MEM[8104] + MEM[8704];
assign MEM[14834] = MEM[8109] + MEM[11370];
assign MEM[14835] = MEM[8124] + MEM[9386];
assign MEM[14836] = MEM[8127] + MEM[9964];
assign MEM[14837] = MEM[8148] + MEM[8854];
assign MEM[14838] = MEM[8159] + MEM[9085];
assign MEM[14839] = MEM[8182] + MEM[8941];
assign MEM[14840] = MEM[8183] + MEM[9627];
assign MEM[14841] = MEM[8184] + MEM[8442];
assign MEM[14842] = MEM[8185] + MEM[9400];
assign MEM[14843] = MEM[8188] + MEM[9665];
assign MEM[14844] = MEM[8189] + MEM[9662];
assign MEM[14845] = MEM[8194] + MEM[8550];
assign MEM[14846] = MEM[8195] + MEM[8419];
assign MEM[14847] = MEM[8200] + MEM[8698];
assign MEM[14848] = MEM[8209] + MEM[8389];
assign MEM[14849] = MEM[8215] + MEM[8631];
assign MEM[14850] = MEM[8229] + MEM[8458];
assign MEM[14851] = MEM[8230] + MEM[8852];
assign MEM[14852] = MEM[8234] + MEM[8379];
assign MEM[14853] = MEM[8248] + MEM[8462];
assign MEM[14854] = MEM[8249] + MEM[8770];
assign MEM[14855] = MEM[8267] + MEM[8575];
assign MEM[14856] = MEM[8271] + MEM[8446];
assign MEM[14857] = MEM[8276] + MEM[5109];
assign MEM[14858] = MEM[8279] + MEM[10055];
assign MEM[14859] = MEM[8281] + MEM[8589];
assign MEM[14860] = MEM[8305] + MEM[11027];
assign MEM[14861] = MEM[8312] + MEM[9136];
assign MEM[14862] = MEM[8313] + MEM[8906];
assign MEM[14863] = MEM[8316] + MEM[10182];
assign MEM[14864] = MEM[8318] + MEM[8439];
assign MEM[14865] = MEM[8321] + MEM[9613];
assign MEM[14866] = MEM[8325] + MEM[9427];
assign MEM[14867] = MEM[8327] + MEM[9050];
assign MEM[14868] = MEM[8329] + MEM[8617];
assign MEM[14869] = MEM[8334] + MEM[8613];
assign MEM[14870] = MEM[8340] + MEM[8649];
assign MEM[14871] = MEM[8346] + MEM[8416];
assign MEM[14872] = MEM[8356] + MEM[2454];
assign MEM[14873] = MEM[8363] + MEM[8881];
assign MEM[14874] = MEM[8367] + MEM[8444];
assign MEM[14875] = MEM[8372] + MEM[11050];
assign MEM[14876] = MEM[8377] + MEM[8530];
assign MEM[14877] = MEM[8378] + MEM[9198];
assign MEM[14878] = MEM[8381] + MEM[8632];
assign MEM[14879] = MEM[8383] + MEM[3150];
assign MEM[14880] = MEM[8385] + MEM[3443];
assign MEM[14881] = MEM[8388] + MEM[8354];
assign MEM[14882] = MEM[8390] + MEM[9122];
assign MEM[14883] = MEM[8392] + MEM[10022];
assign MEM[14884] = MEM[8397] + MEM[9447];
assign MEM[14885] = MEM[8401] + MEM[8694];
assign MEM[14886] = MEM[8402] + MEM[9560];
assign MEM[14887] = MEM[8403] + MEM[8973];
assign MEM[14888] = MEM[8405] + MEM[9352];
assign MEM[14889] = MEM[8406] + MEM[10171];
assign MEM[14890] = MEM[8412] + MEM[8659];
assign MEM[14891] = MEM[8424] + MEM[8619];
assign MEM[14892] = MEM[8436] + MEM[9751];
assign MEM[14893] = MEM[8437] + MEM[8612];
assign MEM[14894] = MEM[8440] + MEM[8787];
assign MEM[14895] = MEM[8441] + MEM[9578];
assign MEM[14896] = MEM[8447] + MEM[10751];
assign MEM[14897] = MEM[8451] + MEM[9318];
assign MEM[14898] = MEM[8452] + MEM[11036];
assign MEM[14899] = MEM[8464] + MEM[9041];
assign MEM[14900] = MEM[8466] + MEM[8889];
assign MEM[14901] = MEM[8478] + MEM[9037];
assign MEM[14902] = MEM[8486] + MEM[8963];
assign MEM[14903] = MEM[8487] + MEM[10083];
assign MEM[14904] = MEM[8491] + MEM[9793];
assign MEM[14905] = MEM[8494] + MEM[9116];
assign MEM[14906] = MEM[8498] + MEM[9096];
assign MEM[14907] = MEM[8499] + MEM[8614];
assign MEM[14908] = MEM[8505] + MEM[9830];
assign MEM[14909] = MEM[8515] + MEM[9152];
assign MEM[14910] = MEM[8517] + MEM[9245];
assign MEM[14911] = MEM[8525] + MEM[9566];
assign MEM[14912] = MEM[8532] + MEM[8988];
assign MEM[14913] = MEM[8534] + MEM[8133];
assign MEM[14914] = MEM[8539] + MEM[9093];
assign MEM[14915] = MEM[8540] + MEM[11188];
assign MEM[14916] = MEM[8542] + MEM[8558];
assign MEM[14917] = MEM[8546] + MEM[9034];
assign MEM[14918] = MEM[8554] + MEM[744];
assign MEM[14919] = MEM[8562] + MEM[8860];
assign MEM[14920] = MEM[8565] + MEM[9180];
assign MEM[14921] = MEM[8567] + MEM[9897];
assign MEM[14922] = MEM[8570] + MEM[4869];
assign MEM[14923] = MEM[8573] + MEM[8949];
assign MEM[14924] = MEM[8574] + MEM[9013];
assign MEM[14925] = MEM[8578] + MEM[3253];
assign MEM[14926] = MEM[8579] + MEM[8712];
assign MEM[14927] = MEM[8588] + MEM[8769];
assign MEM[14928] = MEM[8597] + MEM[8932];
assign MEM[14929] = MEM[8599] + MEM[9780];
assign MEM[14930] = MEM[8600] + MEM[9370];
assign MEM[14931] = MEM[8601] + MEM[10145];
assign MEM[14932] = MEM[8603] + MEM[9795];
assign MEM[14933] = MEM[8611] + MEM[1258];
assign MEM[14934] = MEM[8618] + MEM[9078];
assign MEM[14935] = MEM[8630] + MEM[9553];
assign MEM[14936] = MEM[8637] + MEM[9231];
assign MEM[14937] = MEM[8638] + MEM[9397];
assign MEM[14938] = MEM[8646] + MEM[9211];
assign MEM[14939] = MEM[8647] + MEM[8999];
assign MEM[14940] = MEM[8648] + MEM[9526];
assign MEM[14941] = MEM[8655] + MEM[7706];
assign MEM[14942] = MEM[8660] + MEM[1902];
assign MEM[14943] = MEM[8667] + MEM[8983];
assign MEM[14944] = MEM[8672] + MEM[8795];
assign MEM[14945] = MEM[8677] + MEM[4555];
assign MEM[14946] = MEM[8678] + MEM[10191];
assign MEM[14947] = MEM[8682] + MEM[10265];
assign MEM[14948] = MEM[8686] + MEM[10221];
assign MEM[14949] = MEM[8690] + MEM[8700];
assign MEM[14950] = MEM[8699] + MEM[9254];
assign MEM[14951] = MEM[8707] + MEM[11240];
assign MEM[14952] = MEM[8709] + MEM[11090];
assign MEM[14953] = MEM[8710] + MEM[9794];
assign MEM[14954] = MEM[8711] + MEM[9284];
assign MEM[14955] = MEM[8714] + MEM[9469];
assign MEM[14956] = MEM[8718] + MEM[8952];
assign MEM[14957] = MEM[8719] + MEM[8827];
assign MEM[14958] = MEM[8720] + MEM[7381];
assign MEM[14959] = MEM[8723] + MEM[8410];
assign MEM[14960] = MEM[8728] + MEM[9008];
assign MEM[14961] = MEM[8729] + MEM[10108];
assign MEM[14962] = MEM[8735] + MEM[9423];
assign MEM[14963] = MEM[8750] + MEM[3718];
assign MEM[14964] = MEM[8754] + MEM[9675];
assign MEM[14965] = MEM[8755] + MEM[9572];
assign MEM[14966] = MEM[8760] + MEM[9150];
assign MEM[14967] = MEM[8763] + MEM[8896];
assign MEM[14968] = MEM[8765] + MEM[8981];
assign MEM[14969] = MEM[8766] + MEM[10714];
assign MEM[14970] = MEM[8768] + MEM[9708];
assign MEM[14971] = MEM[8773] + MEM[11325];
assign MEM[14972] = MEM[8774] + MEM[9332];
assign MEM[14973] = MEM[8786] + MEM[11182];
assign MEM[14974] = MEM[8789] + MEM[851];
assign MEM[14975] = MEM[8791] + MEM[10487];
assign MEM[14976] = MEM[8797] + MEM[9200];
assign MEM[14977] = MEM[8806] + MEM[11200];
assign MEM[14978] = MEM[8810] + MEM[9424];
assign MEM[14979] = MEM[8812] + MEM[9885];
assign MEM[14980] = MEM[8820] + MEM[7375];
assign MEM[14981] = MEM[8824] + MEM[9800];
assign MEM[14982] = MEM[8831] + MEM[10958];
assign MEM[14983] = MEM[8833] + MEM[8948];
assign MEM[14984] = MEM[8839] + MEM[9282];
assign MEM[14985] = MEM[8842] + MEM[5895];
assign MEM[14986] = MEM[8843] + MEM[9187];
assign MEM[14987] = MEM[8845] + MEM[9244];
assign MEM[14988] = MEM[8846] + MEM[9260];
assign MEM[14989] = MEM[8847] + MEM[10660];
assign MEM[14990] = MEM[8852] + MEM[10968];
assign MEM[14991] = MEM[8856] + MEM[9411];
assign MEM[14992] = MEM[8858] + MEM[9125];
assign MEM[14993] = MEM[8859] + MEM[9105];
assign MEM[14994] = MEM[8862] + MEM[9262];
assign MEM[14995] = MEM[8871] + MEM[1002];
assign MEM[14996] = MEM[8872] + MEM[9940];
assign MEM[14997] = MEM[8874] + MEM[10864];
assign MEM[14998] = MEM[8877] + MEM[11000];
assign MEM[14999] = MEM[8878] + MEM[11265];
assign MEM[15000] = MEM[8880] + MEM[9887];
assign MEM[15001] = MEM[8882] + MEM[10067];
assign MEM[15002] = MEM[8884] + MEM[11047];
assign MEM[15003] = MEM[8897] + MEM[9529];
assign MEM[15004] = MEM[8898] + MEM[9905];
assign MEM[15005] = MEM[8899] + MEM[10965];
assign MEM[15006] = MEM[8901] + MEM[9435];
assign MEM[15007] = MEM[8903] + MEM[8971];
assign MEM[15008] = MEM[8908] + MEM[10046];
assign MEM[15009] = MEM[8913] + MEM[11306];
assign MEM[15010] = MEM[8919] + MEM[9405];
assign MEM[15011] = MEM[8920] + MEM[9658];
assign MEM[15012] = MEM[8922] + MEM[9002];
assign MEM[15013] = MEM[8926] + MEM[9484];
assign MEM[15014] = MEM[8935] + MEM[10724];
assign MEM[15015] = MEM[8938] + MEM[10338];
assign MEM[15016] = MEM[8945] + MEM[9259];
assign MEM[15017] = MEM[8950] + MEM[10061];
assign MEM[15018] = MEM[8955] + MEM[9237];
assign MEM[15019] = MEM[8956] + MEM[9010];
assign MEM[15020] = MEM[8958] + MEM[11063];
assign MEM[15021] = MEM[8960] + MEM[8936];
assign MEM[15022] = MEM[8968] + MEM[10485];
assign MEM[15023] = MEM[8969] + MEM[10790];
assign MEM[15024] = MEM[8969] + MEM[11057];
assign MEM[15025] = MEM[8982] + MEM[9770];
assign MEM[15026] = MEM[8984] + MEM[10565];
assign MEM[15027] = MEM[8990] + MEM[9615];
assign MEM[15028] = MEM[8996] + MEM[6747];
assign MEM[15029] = MEM[9004] + MEM[10293];
assign MEM[15030] = MEM[9006] + MEM[10281];
assign MEM[15031] = MEM[9011] + MEM[11128];
assign MEM[15032] = MEM[9012] + MEM[9132];
assign MEM[15033] = MEM[9014] + MEM[10930];
assign MEM[15034] = MEM[9017] + MEM[7125];
assign MEM[15035] = MEM[9021] + MEM[9049];
assign MEM[15036] = MEM[9023] + MEM[9577];
assign MEM[15037] = MEM[9024] + MEM[9380];
assign MEM[15038] = MEM[9027] + MEM[9541];
assign MEM[15039] = MEM[9030] + MEM[9573];
assign MEM[15040] = MEM[9032] + MEM[9248];
assign MEM[15041] = MEM[9033] + MEM[9786];
assign MEM[15042] = MEM[9038] + MEM[9372];
assign MEM[15043] = MEM[9047] + MEM[10172];
assign MEM[15044] = MEM[9056] + MEM[9222];
assign MEM[15045] = MEM[9058] + MEM[10415];
assign MEM[15046] = MEM[9063] + MEM[9206];
assign MEM[15047] = MEM[9066] + MEM[10052];
assign MEM[15048] = MEM[9069] + MEM[9339];
assign MEM[15049] = MEM[9070] + MEM[11796];
assign MEM[15050] = MEM[9072] + MEM[9288];
assign MEM[15051] = MEM[9073] + MEM[11004];
assign MEM[15052] = MEM[9074] + MEM[10054];
assign MEM[15053] = MEM[9074] + MEM[11115];
assign MEM[15054] = MEM[9075] + MEM[9440];
assign MEM[15055] = MEM[9076] + MEM[11016];
assign MEM[15056] = MEM[9079] + MEM[8140];
assign MEM[15057] = MEM[9082] + MEM[10863];
assign MEM[15058] = MEM[9084] + MEM[9820];
assign MEM[15059] = MEM[9095] + MEM[11119];
assign MEM[15060] = MEM[9097] + MEM[9174];
assign MEM[15061] = MEM[9098] + MEM[9133];
assign MEM[15062] = MEM[9100] + MEM[9503];
assign MEM[15063] = MEM[9108] + MEM[10081];
assign MEM[15064] = MEM[9111] + MEM[9849];
assign MEM[15065] = MEM[9112] + MEM[9343];
assign MEM[15066] = MEM[9115] + MEM[9518];
assign MEM[15067] = MEM[9118] + MEM[9363];
assign MEM[15068] = MEM[9121] + MEM[9141];
assign MEM[15069] = MEM[9123] + MEM[9345];
assign MEM[15070] = MEM[9124] + MEM[11317];
assign MEM[15071] = MEM[9128] + MEM[10311];
assign MEM[15072] = MEM[9129] + MEM[9457];
assign MEM[15073] = MEM[9131] + MEM[9985];
assign MEM[15074] = MEM[9134] + MEM[9874];
assign MEM[15075] = MEM[9138] + MEM[10949];
assign MEM[15076] = MEM[9140] + MEM[9668];
assign MEM[15077] = MEM[9144] + MEM[10279];
assign MEM[15078] = MEM[9146] + MEM[8177];
assign MEM[15079] = MEM[9151] + MEM[10077];
assign MEM[15080] = MEM[9165] + MEM[9596];
assign MEM[15081] = MEM[9172] + MEM[10806];
assign MEM[15082] = MEM[9176] + MEM[10912];
assign MEM[15083] = MEM[9189] + MEM[9519];
assign MEM[15084] = MEM[9194] + MEM[10312];
assign MEM[15085] = MEM[9196] + MEM[11006];
assign MEM[15086] = MEM[9197] + MEM[9642];
assign MEM[15087] = MEM[9202] + MEM[9501];
assign MEM[15088] = MEM[9205] + MEM[810];
assign MEM[15089] = MEM[9209] + MEM[9342];
assign MEM[15090] = MEM[9210] + MEM[10217];
assign MEM[15091] = MEM[9212] + MEM[10923];
assign MEM[15092] = MEM[9224] + MEM[10031];
assign MEM[15093] = MEM[9243] + MEM[1643];
assign MEM[15094] = MEM[9246] + MEM[9479];
assign MEM[15095] = MEM[9249] + MEM[11024];
assign MEM[15096] = MEM[9250] + MEM[10039];
assign MEM[15097] = MEM[9252] + MEM[9310];
assign MEM[15098] = MEM[9266] + MEM[9720];
assign MEM[15099] = MEM[9267] + MEM[11509];
assign MEM[15100] = MEM[9270] + MEM[11201];
assign MEM[15101] = MEM[9273] + MEM[9239];
assign MEM[15102] = MEM[9277] + MEM[9845];
assign MEM[15103] = MEM[9281] + MEM[9359];
assign MEM[15104] = MEM[9282] + MEM[11236];
assign MEM[15105] = MEM[9294] + MEM[9590];
assign MEM[15106] = MEM[9300] + MEM[9344];
assign MEM[15107] = MEM[9301] + MEM[9500];
assign MEM[15108] = MEM[9305] + MEM[9836];
assign MEM[15109] = MEM[9312] + MEM[9381];
assign MEM[15110] = MEM[9319] + MEM[9341];
assign MEM[15111] = MEM[9321] + MEM[9729];
assign MEM[15112] = MEM[9323] + MEM[10176];
assign MEM[15113] = MEM[9325] + MEM[10246];
assign MEM[15114] = MEM[9326] + MEM[9696];
assign MEM[15115] = MEM[9328] + MEM[9495];
assign MEM[15116] = MEM[9329] + MEM[9595];
assign MEM[15117] = MEM[9333] + MEM[11029];
assign MEM[15118] = MEM[9336] + MEM[11058];
assign MEM[15119] = MEM[9340] + MEM[9369];
assign MEM[15120] = MEM[9346] + MEM[9682];
assign MEM[15121] = MEM[9348] + MEM[11126];
assign MEM[15122] = MEM[9351] + MEM[9474];
assign MEM[15123] = MEM[9358] + MEM[9364];
assign MEM[15124] = MEM[9362] + MEM[10260];
assign MEM[15125] = MEM[9365] + MEM[9635];
assign MEM[15126] = MEM[9377] + MEM[11464];
assign MEM[15127] = MEM[9382] + MEM[10096];
assign MEM[15128] = MEM[9385] + MEM[10100];
assign MEM[15129] = MEM[9393] + MEM[9601];
assign MEM[15130] = MEM[9395] + MEM[10131];
assign MEM[15131] = MEM[9401] + MEM[9813];
assign MEM[15132] = MEM[9402] + MEM[10110];
assign MEM[15133] = MEM[9404] + MEM[9678];
assign MEM[15134] = MEM[9412] + MEM[9317];
assign MEM[15135] = MEM[9413] + MEM[10383];
assign MEM[15136] = MEM[9414] + MEM[10027];
assign MEM[15137] = MEM[9418] + MEM[10124];
assign MEM[15138] = MEM[9421] + MEM[11198];
assign MEM[15139] = MEM[9425] + MEM[9016];
assign MEM[15140] = MEM[9432] + MEM[11062];
assign MEM[15141] = MEM[9434] + MEM[11139];
assign MEM[15142] = MEM[9436] + MEM[9594];
assign MEM[15143] = MEM[9439] + MEM[8580];
assign MEM[15144] = MEM[9442] + MEM[9552];
assign MEM[15145] = MEM[9444] + MEM[10090];
assign MEM[15146] = MEM[9452] + MEM[9064];
assign MEM[15147] = MEM[9456] + MEM[11065];
assign MEM[15148] = MEM[9459] + MEM[10232];
assign MEM[15149] = MEM[9462] + MEM[7071];
assign MEM[15150] = MEM[9470] + MEM[11124];
assign MEM[15151] = MEM[9471] + MEM[8904];
assign MEM[15152] = MEM[9473] + MEM[9785];
assign MEM[15153] = MEM[9475] + MEM[10051];
assign MEM[15154] = MEM[9477] + MEM[9697];
assign MEM[15155] = MEM[9482] + MEM[10036];
assign MEM[15156] = MEM[9491] + MEM[11014];
assign MEM[15157] = MEM[9492] + MEM[9598];
assign MEM[15158] = MEM[9493] + MEM[9545];
assign MEM[15159] = MEM[9496] + MEM[9761];
assign MEM[15160] = MEM[9497] + MEM[10642];
assign MEM[15161] = MEM[9498] + MEM[10966];
assign MEM[15162] = MEM[9509] + MEM[10183];
assign MEM[15163] = MEM[9512] + MEM[11129];
assign MEM[15164] = MEM[9517] + MEM[562];
assign MEM[15165] = MEM[9520] + MEM[9666];
assign MEM[15166] = MEM[9534] + MEM[11031];
assign MEM[15167] = MEM[9536] + MEM[10983];
assign MEM[15168] = MEM[9548] + MEM[9722];
assign MEM[15169] = MEM[9556] + MEM[10817];
assign MEM[15170] = MEM[9559] + MEM[8972];
assign MEM[15171] = MEM[9561] + MEM[10139];
assign MEM[15172] = MEM[9575] + MEM[10376];
assign MEM[15173] = MEM[9579] + MEM[10980];
assign MEM[15174] = MEM[9582] + MEM[9863];
assign MEM[15175] = MEM[9592] + MEM[9963];
assign MEM[15176] = MEM[9603] + MEM[10474];
assign MEM[15177] = MEM[9605] + MEM[9797];
assign MEM[15178] = MEM[9608] + MEM[10943];
assign MEM[15179] = MEM[9609] + MEM[7775];
assign MEM[15180] = MEM[9610] + MEM[8970];
assign MEM[15181] = MEM[9611] + MEM[11053];
assign MEM[15182] = MEM[9622] + MEM[10076];
assign MEM[15183] = MEM[9623] + MEM[8431];
assign MEM[15184] = MEM[9626] + MEM[11048];
assign MEM[15185] = MEM[9628] + MEM[10148];
assign MEM[15186] = MEM[9629] + MEM[7460];
assign MEM[15187] = MEM[9630] + MEM[10566];
assign MEM[15188] = MEM[9634] + MEM[11484];
assign MEM[15189] = MEM[9639] + MEM[6956];
assign MEM[15190] = MEM[9644] + MEM[10168];
assign MEM[15191] = MEM[9645] + MEM[10963];
assign MEM[15192] = MEM[9647] + MEM[11261];
assign MEM[15193] = MEM[9654] + MEM[9882];
assign MEM[15194] = MEM[9657] + MEM[11059];
assign MEM[15195] = MEM[9660] + MEM[9856];
assign MEM[15196] = MEM[9661] + MEM[9923];
assign MEM[15197] = MEM[9670] + MEM[11100];
assign MEM[15198] = MEM[9679] + MEM[10078];
assign MEM[15199] = MEM[9680] + MEM[11061];
assign MEM[15200] = MEM[9686] + MEM[10121];
assign MEM[15201] = MEM[9687] + MEM[10894];
assign MEM[15202] = MEM[9689] + MEM[10879];
assign MEM[15203] = MEM[9690] + MEM[9417];
assign MEM[15204] = MEM[9704] + MEM[9747];
assign MEM[15205] = MEM[9710] + MEM[11271];
assign MEM[15206] = MEM[9715] + MEM[11143];
assign MEM[15207] = MEM[9719] + MEM[7286];
assign MEM[15208] = MEM[9731] + MEM[10038];
assign MEM[15209] = MEM[9732] + MEM[10005];
assign MEM[15210] = MEM[9738] + MEM[11148];
assign MEM[15211] = MEM[9740] + MEM[9829];
assign MEM[15212] = MEM[9752] + MEM[11067];
assign MEM[15213] = MEM[9756] + MEM[10742];
assign MEM[15214] = MEM[9759] + MEM[10667];
assign MEM[15215] = MEM[9764] + MEM[10879];
assign MEM[15216] = MEM[9768] + MEM[11083];
assign MEM[15217] = MEM[9776] + MEM[9408];
assign MEM[15218] = MEM[9787] + MEM[9945];
assign MEM[15219] = MEM[9789] + MEM[11605];
assign MEM[15220] = MEM[9799] + MEM[9916];
assign MEM[15221] = MEM[9809] + MEM[9828];
assign MEM[15222] = MEM[9819] + MEM[9168];
assign MEM[15223] = MEM[9823] + MEM[5508];
assign MEM[15224] = MEM[9824] + MEM[11051];
assign MEM[15225] = MEM[9825] + MEM[9918];
assign MEM[15226] = MEM[9842] + MEM[10041];
assign MEM[15227] = MEM[9843] + MEM[10354];
assign MEM[15228] = MEM[9864] + MEM[11380];
assign MEM[15229] = MEM[9890] + MEM[11331];
assign MEM[15230] = MEM[9901] + MEM[10141];
assign MEM[15231] = MEM[9911] + MEM[11324];
assign MEM[15232] = MEM[9915] + MEM[9909];
assign MEM[15233] = MEM[9919] + MEM[754];
assign MEM[15234] = MEM[9924] + MEM[9854];
assign MEM[15235] = MEM[9927] + MEM[11141];
assign MEM[15236] = MEM[9933] + MEM[10018];
assign MEM[15237] = MEM[9934] + MEM[9304];
assign MEM[15238] = MEM[9941] + MEM[9298];
assign MEM[15239] = MEM[9944] + MEM[10989];
assign MEM[15240] = MEM[9947] + MEM[10569];
assign MEM[15241] = MEM[9952] + MEM[10364];
assign MEM[15242] = MEM[9956] + MEM[9943];
assign MEM[15243] = MEM[9958] + MEM[10913];
assign MEM[15244] = MEM[9968] + MEM[10136];
assign MEM[15245] = MEM[9972] + MEM[9685];
assign MEM[15246] = MEM[9973] + MEM[10912];
assign MEM[15247] = MEM[9974] + MEM[10955];
assign MEM[15248] = MEM[9976] + MEM[10114];
assign MEM[15249] = MEM[9982] + MEM[10901];
assign MEM[15250] = MEM[9984] + MEM[6723];
assign MEM[15251] = MEM[9989] + MEM[8779];
assign MEM[15252] = MEM[9992] + MEM[11423];
assign MEM[15253] = MEM[10000] + MEM[10783];
assign MEM[15254] = MEM[10002] + MEM[10382];
assign MEM[15255] = MEM[10011] + MEM[5429];
assign MEM[15256] = MEM[10015] + MEM[9816];
assign MEM[15257] = MEM[10023] + MEM[10044];
assign MEM[15258] = MEM[10047] + MEM[11191];
assign MEM[15259] = MEM[10049] + MEM[9962];
assign MEM[15260] = MEM[10071] + MEM[10979];
assign MEM[15261] = MEM[10080] + MEM[11160];
assign MEM[15262] = MEM[10085] + MEM[4187];
assign MEM[15263] = MEM[10091] + MEM[10060];
assign MEM[15264] = MEM[10094] + MEM[9749];
assign MEM[15265] = MEM[10095] + MEM[12424];
assign MEM[15266] = MEM[10116] + MEM[10098];
assign MEM[15267] = MEM[10129] + MEM[9993];
assign MEM[15268] = MEM[10164] + MEM[11118];
assign MEM[15269] = MEM[10177] + MEM[10305];
assign MEM[15270] = MEM[10194] + MEM[5078];
assign MEM[15271] = MEM[10203] + MEM[11013];
assign MEM[15272] = MEM[10212] + MEM[12240];
assign MEM[15273] = MEM[10216] + MEM[2739];
assign MEM[15274] = MEM[10218] + MEM[10045];
assign MEM[15275] = MEM[10223] + MEM[11035];
assign MEM[15276] = MEM[10245] + MEM[2806];
assign MEM[15277] = MEM[10249] + MEM[11146];
assign MEM[15278] = MEM[10250] + MEM[10914];
assign MEM[15279] = MEM[10251] + MEM[11427];
assign MEM[15280] = MEM[10262] + MEM[11844];
assign MEM[15281] = MEM[10288] + MEM[10921];
assign MEM[15282] = MEM[10325] + MEM[9003];
assign MEM[15283] = MEM[10327] + MEM[11298];
assign MEM[15284] = MEM[10335] + MEM[2542];
assign MEM[15285] = MEM[10340] + MEM[11589];
assign MEM[15286] = MEM[10345] + MEM[11078];
assign MEM[15287] = MEM[10351] + MEM[10257];
assign MEM[15288] = MEM[10356] + MEM[11049];
assign MEM[15289] = MEM[10369] + MEM[3655];
assign MEM[15290] = MEM[10386] + MEM[990];
assign MEM[15291] = MEM[10390] + MEM[11070];
assign MEM[15292] = MEM[10391] + MEM[10406];
assign MEM[15293] = MEM[10426] + MEM[10437];
assign MEM[15294] = MEM[10456] + MEM[9420];
assign MEM[15295] = MEM[10527] + MEM[10444];
assign MEM[15296] = MEM[10535] + MEM[11798];
assign MEM[15297] = MEM[10635] + MEM[10972];
assign MEM[15298] = MEM[10666] + MEM[11172];
assign MEM[15299] = MEM[10710] + MEM[10975];
assign MEM[15300] = MEM[10715] + MEM[12248];
assign MEM[15301] = MEM[10760] + MEM[10925];
assign MEM[15302] = MEM[10822] + MEM[4123];
assign MEM[15303] = MEM[10880] + MEM[11246];
assign MEM[15304] = MEM[10888] + MEM[6444];
assign MEM[15305] = MEM[10889] + MEM[10301];
assign MEM[15306] = MEM[10890] + MEM[10329];
assign MEM[15307] = MEM[10892] + MEM[9335];
assign MEM[15308] = MEM[10907] + MEM[11189];
assign MEM[15309] = MEM[10915] + MEM[7856];
assign MEM[15310] = MEM[10920] + MEM[8943];
assign MEM[15311] = MEM[10932] + MEM[6014];
assign MEM[15312] = MEM[10933] + MEM[1846];
assign MEM[15313] = MEM[10939] + MEM[10404];
assign MEM[15314] = MEM[10942] + MEM[10875];
assign MEM[15315] = MEM[10944] + MEM[9925];
assign MEM[15316] = MEM[10953] + MEM[10237];
assign MEM[15317] = MEM[10957] + MEM[6206];
assign MEM[15318] = MEM[10961] + MEM[9881];
assign MEM[15319] = MEM[10977] + MEM[8541];
assign MEM[15320] = MEM[10987] + MEM[10313];
assign MEM[15321] = MEM[10990] + MEM[12672];
assign MEM[15322] = MEM[10991] + MEM[9036];
assign MEM[15323] = MEM[10992] + MEM[7070];
assign MEM[15324] = MEM[11002] + MEM[10555];
assign MEM[15325] = MEM[11009] + MEM[10374];
assign MEM[15326] = MEM[11015] + MEM[11319];
assign MEM[15327] = MEM[11018] + MEM[9221];
assign MEM[15328] = MEM[11028] + MEM[11264];
assign MEM[15329] = MEM[11033] + MEM[858];
assign MEM[15330] = MEM[11034] + MEM[11158];
assign MEM[15331] = MEM[11037] + MEM[1284];
assign MEM[15332] = MEM[11040] + MEM[10062];
assign MEM[15333] = MEM[11041] + MEM[9938];
assign MEM[15334] = MEM[11042] + MEM[8931];
assign MEM[15335] = MEM[11045] + MEM[11543];
assign MEM[15336] = MEM[11046] + MEM[11109];
assign MEM[15337] = MEM[11052] + MEM[11250];
assign MEM[15338] = MEM[11055] + MEM[1366];
assign MEM[15339] = MEM[11056] + MEM[6939];
assign MEM[15340] = MEM[11060] + MEM[9147];
assign MEM[15341] = MEM[11066] + MEM[9818];
assign MEM[15342] = MEM[11069] + MEM[11002];
assign MEM[15343] = MEM[11073] + MEM[10503];
assign MEM[15344] = MEM[11073] + MEM[11665];
assign MEM[15345] = MEM[11074] + MEM[3442];
assign MEM[15346] = MEM[11075] + MEM[11357];
assign MEM[15347] = MEM[11076] + MEM[9516];
assign MEM[15348] = MEM[11077] + MEM[10530];
assign MEM[15349] = MEM[11079] + MEM[3178];
assign MEM[15350] = MEM[11080] + MEM[9502];
assign MEM[15351] = MEM[11082] + MEM[10702];
assign MEM[15352] = MEM[11082] + MEM[11252];
assign MEM[15353] = MEM[11085] + MEM[9521];
assign MEM[15354] = MEM[11088] + MEM[11341];
assign MEM[15355] = MEM[11091] + MEM[11137];
assign MEM[15356] = MEM[11094] + MEM[9815];
assign MEM[15357] = MEM[11096] + MEM[11322];
assign MEM[15358] = MEM[11098] + MEM[11199];
assign MEM[15359] = MEM[11103] + MEM[9677];
assign MEM[15360] = MEM[11106] + MEM[11110];
assign MEM[15361] = MEM[11112] + MEM[10475];
assign MEM[15362] = MEM[11113] + MEM[11142];
assign MEM[15363] = MEM[11114] + MEM[9407];
assign MEM[15364] = MEM[11123] + MEM[5571];
assign MEM[15365] = MEM[11125] + MEM[11194];
assign MEM[15366] = MEM[11127] + MEM[10945];
assign MEM[15367] = MEM[11130] + MEM[11136];
assign MEM[15368] = MEM[11134] + MEM[11168];
assign MEM[15369] = MEM[11135] + MEM[9694];
assign MEM[15370] = MEM[11140] + MEM[9307];
assign MEM[15371] = MEM[11144] + MEM[9655];
assign MEM[15372] = MEM[11145] + MEM[9953];
assign MEM[15373] = MEM[11147] + MEM[5986];
assign MEM[15374] = MEM[11149] + MEM[4885];
assign MEM[15375] = MEM[11152] + MEM[11245];
assign MEM[15376] = MEM[11153] + MEM[8918];
assign MEM[15377] = MEM[11154] + MEM[11164];
assign MEM[15378] = MEM[11156] + MEM[10206];
assign MEM[15379] = MEM[11156] + MEM[10128];
assign MEM[15380] = MEM[11157] + MEM[11180];
assign MEM[15381] = MEM[11159] + MEM[10596];
assign MEM[15382] = MEM[11162] + MEM[10331];
assign MEM[15383] = MEM[11165] + MEM[11227];
assign MEM[15384] = MEM[11166] + MEM[3555];
assign MEM[15385] = MEM[11167] + MEM[9602];
assign MEM[15386] = MEM[11173] + MEM[10082];
assign MEM[15387] = MEM[11175] + MEM[11411];
assign MEM[15388] = MEM[11176] + MEM[10271];
assign MEM[15389] = MEM[11177] + MEM[9621];
assign MEM[15390] = MEM[11202] + MEM[10558];
assign MEM[15391] = MEM[11205] + MEM[11230];
assign MEM[15392] = MEM[11207] + MEM[9878];
assign MEM[15393] = MEM[11209] + MEM[11501];
assign MEM[15394] = MEM[11211] + MEM[11150];
assign MEM[15395] = MEM[11219] + MEM[10344];
assign MEM[15396] = MEM[11224] + MEM[7963];
assign MEM[15397] = MEM[11235] + MEM[8269];
assign MEM[15398] = MEM[11242] + MEM[8475];
assign MEM[15399] = MEM[11243] + MEM[10465];
assign MEM[15400] = MEM[11247] + MEM[3413];
assign MEM[15401] = MEM[11257] + MEM[11919];
assign MEM[15402] = MEM[11259] + MEM[11260];
assign MEM[15403] = MEM[11262] + MEM[11395];
assign MEM[15404] = MEM[11267] + MEM[13469];
assign MEM[15405] = MEM[11269] + MEM[9562];
assign MEM[15406] = MEM[11270] + MEM[11305];
assign MEM[15407] = MEM[11272] + MEM[11348];
assign MEM[15408] = MEM[11275] + MEM[9955];
assign MEM[15409] = MEM[11283] + MEM[11332];
assign MEM[15410] = MEM[11285] + MEM[11935];
assign MEM[15411] = MEM[11286] + MEM[11473];
assign MEM[15412] = MEM[11289] + MEM[10079];
assign MEM[15413] = MEM[11296] + MEM[5124];
assign MEM[15414] = MEM[11297] + MEM[10774];
assign MEM[15415] = MEM[11313] + MEM[11383];
assign MEM[15416] = MEM[11315] + MEM[3526];
assign MEM[15417] = MEM[11316] + MEM[9489];
assign MEM[15418] = MEM[11330] + MEM[1259];
assign MEM[15419] = MEM[11334] + MEM[11849];
assign MEM[15420] = MEM[11369] + MEM[13025];
assign MEM[15421] = MEM[11391] + MEM[11206];
assign MEM[15422] = MEM[11403] + MEM[8193];
assign MEM[15423] = MEM[11408] + MEM[11806];
assign MEM[15424] = MEM[11440] + MEM[7916];
assign MEM[15425] = MEM[11445] + MEM[4799];
assign MEM[15426] = MEM[11447] + MEM[11095];
assign MEM[15427] = MEM[11459] + MEM[11502];
assign MEM[15428] = MEM[11477] + MEM[4677];
assign MEM[15429] = MEM[11478] + MEM[9807];
assign MEM[15430] = MEM[11490] + MEM[10034];
assign MEM[15431] = MEM[11516] + MEM[11338];
assign MEM[15432] = MEM[11524] + MEM[10225];
assign MEM[15433] = MEM[11526] + MEM[8456];
assign MEM[15434] = MEM[11550] + MEM[10733];
assign MEM[15435] = MEM[11558] + MEM[4627];
assign MEM[15436] = MEM[11652] + MEM[10029];
assign MEM[15437] = MEM[11741] + MEM[9524];
assign MEM[15438] = MEM[11795] + MEM[8725];
assign MEM[15439] = MEM[11864] + MEM[9255];
assign MEM[15440] = MEM[11873] + MEM[9880];
assign MEM[15441] = MEM[11889] + MEM[11020];
assign MEM[15442] = MEM[13111] + MEM[11033];
assign MEM[15443] = MEM[13874] + MEM[8781];
assign MEM[15444] = MEM[14097] + MEM[11973];
assign MEM[15445] = MEM[14259] + MEM[9110];
assign MEM[15446] = MEM[14287] + MEM[11268];
assign MEM[15447] = MEM[14308] + MEM[9261];
assign MEM[15448] = MEM[14399] + MEM[13453];
assign MEM[15449] = MEM[14870] + MEM[9303];
assign MEM[15450] = MEM[15407] + MEM[11848];
assign MEM[15451] = MEM[14] + MEM[13263];
assign MEM[15452] = MEM[29] + MEM[13135];
assign MEM[15453] = MEM[37] + MEM[13983];
assign MEM[15454] = MEM[47] + MEM[7279];
assign MEM[15455] = MEM[77] + MEM[13096];
assign MEM[15456] = MEM[85] + MEM[628];
assign MEM[15457] = MEM[101] + MEM[13011];
assign MEM[15458] = MEM[102] + MEM[11452];
assign MEM[15459] = MEM[103] + MEM[10186];
assign MEM[15460] = MEM[111] + MEM[7793];
assign MEM[15461] = MEM[119] + MEM[967];
assign MEM[15462] = MEM[126] + MEM[13411];
assign MEM[15463] = MEM[143] + MEM[1069];
assign MEM[15464] = MEM[189] + MEM[9805];
assign MEM[15465] = MEM[239] + MEM[7146];
assign MEM[15466] = MEM[245] + MEM[9895];
assign MEM[15467] = MEM[246] + MEM[13446];
assign MEM[15468] = MEM[253] + MEM[7817];
assign MEM[15469] = MEM[271] + MEM[11203];
assign MEM[15470] = MEM[291] + MEM[8756];
assign MEM[15471] = MEM[299] + MEM[12507];
assign MEM[15472] = MEM[308] + MEM[7449];
assign MEM[15473] = MEM[334] + MEM[846];
assign MEM[15474] = MEM[346] + MEM[9778];
assign MEM[15475] = MEM[348] + MEM[2963];
assign MEM[15476] = MEM[358] + MEM[9169];
assign MEM[15477] = MEM[362] + MEM[10088];
assign MEM[15478] = MEM[367] + MEM[3038];
assign MEM[15479] = MEM[373] + MEM[6802];
assign MEM[15480] = MEM[375] + MEM[959];
assign MEM[15481] = MEM[386] + MEM[11004];
assign MEM[15482] = MEM[387] + MEM[3557];
assign MEM[15483] = MEM[396] + MEM[7103];
assign MEM[15484] = MEM[397] + MEM[10241];
assign MEM[15485] = MEM[412] + MEM[10458];
assign MEM[15486] = MEM[421] + MEM[7770];
assign MEM[15487] = MEM[430] + MEM[10407];
assign MEM[15488] = MEM[447] + MEM[9773];
assign MEM[15489] = MEM[454] + MEM[11279];
assign MEM[15490] = MEM[462] + MEM[8584];
assign MEM[15491] = MEM[478] + MEM[10278];
assign MEM[15492] = MEM[499] + MEM[2380];
assign MEM[15493] = MEM[500] + MEM[1053];
assign MEM[15494] = MEM[514] + MEM[7258];
assign MEM[15495] = MEM[527] + MEM[2323];
assign MEM[15496] = MEM[530] + MEM[5929];
assign MEM[15497] = MEM[532] + MEM[9865];
assign MEM[15498] = MEM[535] + MEM[11101];
assign MEM[15499] = MEM[538] + MEM[13351];
assign MEM[15500] = MEM[546] + MEM[3238];
assign MEM[15501] = MEM[551] + MEM[11314];
assign MEM[15502] = MEM[578] + MEM[12352];
assign MEM[15503] = MEM[583] + MEM[1012];
assign MEM[15504] = MEM[594] + MEM[8861];
assign MEM[15505] = MEM[597] + MEM[4014];
assign MEM[15506] = MEM[600] + MEM[11299];
assign MEM[15507] = MEM[618] + MEM[7826];
assign MEM[15508] = MEM[621] + MEM[10751];
assign MEM[15509] = MEM[629] + MEM[12451];
assign MEM[15510] = MEM[631] + MEM[8980];
assign MEM[15511] = MEM[646] + MEM[11748];
assign MEM[15512] = MEM[652] + MEM[5581];
assign MEM[15513] = MEM[687] + MEM[12841];
assign MEM[15514] = MEM[701] + MEM[12065];
assign MEM[15515] = MEM[703] + MEM[10657];
assign MEM[15516] = MEM[715] + MEM[7842];
assign MEM[15517] = MEM[718] + MEM[3084];
assign MEM[15518] = MEM[722] + MEM[11487];
assign MEM[15519] = MEM[723] + MEM[9555];
assign MEM[15520] = MEM[727] + MEM[10215];
assign MEM[15521] = MEM[730] + MEM[4374];
assign MEM[15522] = MEM[733] + MEM[7531];
assign MEM[15523] = MEM[743] + MEM[11497];
assign MEM[15524] = MEM[755] + MEM[5285];
assign MEM[15525] = MEM[759] + MEM[9620];
assign MEM[15526] = MEM[772] + MEM[9961];
assign MEM[15527] = MEM[774] + MEM[11517];
assign MEM[15528] = MEM[796] + MEM[9208];
assign MEM[15529] = MEM[804] + MEM[13590];
assign MEM[15530] = MEM[811] + MEM[8684];
assign MEM[15531] = MEM[821] + MEM[10380];
assign MEM[15532] = MEM[835] + MEM[5546];
assign MEM[15533] = MEM[836] + MEM[11434];
assign MEM[15534] = MEM[837] + MEM[9349];
assign MEM[15535] = MEM[838] + MEM[12634];
assign MEM[15536] = MEM[842] + MEM[9892];
assign MEM[15537] = MEM[843] + MEM[10230];
assign MEM[15538] = MEM[850] + MEM[7237];
assign MEM[15539] = MEM[866] + MEM[3867];
assign MEM[15540] = MEM[875] + MEM[7786];
assign MEM[15541] = MEM[887] + MEM[4135];
assign MEM[15542] = MEM[894] + MEM[1100];
assign MEM[15543] = MEM[915] + MEM[4211];
assign MEM[15544] = MEM[917] + MEM[7837];
assign MEM[15545] = MEM[973] + MEM[10270];
assign MEM[15546] = MEM[980] + MEM[2133];
assign MEM[15547] = MEM[982] + MEM[11492];
assign MEM[15548] = MEM[997] + MEM[9192];
assign MEM[15549] = MEM[1003] + MEM[1812];
assign MEM[15550] = MEM[1006] + MEM[7767];
assign MEM[15551] = MEM[1010] + MEM[9990];
assign MEM[15552] = MEM[1036] + MEM[1565];
assign MEM[15553] = MEM[1042] + MEM[8921];
assign MEM[15554] = MEM[1052] + MEM[9394];
assign MEM[15555] = MEM[1066] + MEM[12140];
assign MEM[15556] = MEM[1070] + MEM[6994];
assign MEM[15557] = MEM[1075] + MEM[6972];
assign MEM[15558] = MEM[1077] + MEM[10302];
assign MEM[15559] = MEM[1083] + MEM[9563];
assign MEM[15560] = MEM[1084] + MEM[11455];
assign MEM[15561] = MEM[1087] + MEM[11307];
assign MEM[15562] = MEM[1091] + MEM[9688];
assign MEM[15563] = MEM[1098] + MEM[10616];
assign MEM[15564] = MEM[1117] + MEM[10501];
assign MEM[15565] = MEM[1118] + MEM[14215];
assign MEM[15566] = MEM[1159] + MEM[3658];
assign MEM[15567] = MEM[1163] + MEM[9513];
assign MEM[15568] = MEM[1174] + MEM[7386];
assign MEM[15569] = MEM[1180] + MEM[13399];
assign MEM[15570] = MEM[1181] + MEM[10258];
assign MEM[15571] = MEM[1187] + MEM[9779];
assign MEM[15572] = MEM[1188] + MEM[9977];
assign MEM[15573] = MEM[1198] + MEM[11105];
assign MEM[15574] = MEM[1221] + MEM[9490];
assign MEM[15575] = MEM[1222] + MEM[13207];
assign MEM[15576] = MEM[1231] + MEM[13524];
assign MEM[15577] = MEM[1237] + MEM[11750];
assign MEM[15578] = MEM[1244] + MEM[1823];
assign MEM[15579] = MEM[1245] + MEM[10012];
assign MEM[15580] = MEM[1267] + MEM[11371];
assign MEM[15581] = MEM[1290] + MEM[11468];
assign MEM[15582] = MEM[1301] + MEM[11394];
assign MEM[15583] = MEM[1316] + MEM[10057];
assign MEM[15584] = MEM[1330] + MEM[5797];
assign MEM[15585] = MEM[1333] + MEM[9195];
assign MEM[15586] = MEM[1334] + MEM[13360];
assign MEM[15587] = MEM[1343] + MEM[7887];
assign MEM[15588] = MEM[1365] + MEM[7274];
assign MEM[15589] = MEM[1379] + MEM[7259];
assign MEM[15590] = MEM[1383] + MEM[8514];
assign MEM[15591] = MEM[1391] + MEM[11288];
assign MEM[15592] = MEM[1406] + MEM[6844];
assign MEM[15593] = MEM[1411] + MEM[10348];
assign MEM[15594] = MEM[1412] + MEM[11163];
assign MEM[15595] = MEM[1413] + MEM[11015];
assign MEM[15596] = MEM[1420] + MEM[11100];
assign MEM[15597] = MEM[1431] + MEM[3986];
assign MEM[15598] = MEM[1450] + MEM[3962];
assign MEM[15599] = MEM[1454] + MEM[6992];
assign MEM[15600] = MEM[1459] + MEM[3004];
assign MEM[15601] = MEM[1460] + MEM[11190];
assign MEM[15602] = MEM[1461] + MEM[2245];
assign MEM[15603] = MEM[1466] + MEM[3163];
assign MEM[15604] = MEM[1468] + MEM[10709];
assign MEM[15605] = MEM[1475] + MEM[10155];
assign MEM[15606] = MEM[1482] + MEM[11320];
assign MEM[15607] = MEM[1484] + MEM[12716];
assign MEM[15608] = MEM[1490] + MEM[11746];
assign MEM[15609] = MEM[1493] + MEM[12539];
assign MEM[15610] = MEM[1495] + MEM[8451];
assign MEM[15611] = MEM[1502] + MEM[10987];
assign MEM[15612] = MEM[1524] + MEM[10359];
assign MEM[15613] = MEM[1526] + MEM[10213];
assign MEM[15614] = MEM[1530] + MEM[11996];
assign MEM[15615] = MEM[1533] + MEM[2130];
assign MEM[15616] = MEM[1538] + MEM[2750];
assign MEM[15617] = MEM[1539] + MEM[11238];
assign MEM[15618] = MEM[1541] + MEM[10574];
assign MEM[15619] = MEM[1557] + MEM[9891];
assign MEM[15620] = MEM[1559] + MEM[2630];
assign MEM[15621] = MEM[1567] + MEM[4142];
assign MEM[15622] = MEM[1580] + MEM[7160];
assign MEM[15623] = MEM[1595] + MEM[10065];
assign MEM[15624] = MEM[1603] + MEM[9139];
assign MEM[15625] = MEM[1606] + MEM[12392];
assign MEM[15626] = MEM[1615] + MEM[13505];
assign MEM[15627] = MEM[1618] + MEM[6498];
assign MEM[15628] = MEM[1620] + MEM[11071];
assign MEM[15629] = MEM[1622] + MEM[8288];
assign MEM[15630] = MEM[1631] + MEM[10384];
assign MEM[15631] = MEM[1637] + MEM[12923];
assign MEM[15632] = MEM[1642] + MEM[2653];
assign MEM[15633] = MEM[1642] + MEM[9214];
assign MEM[15634] = MEM[1662] + MEM[8848];
assign MEM[15635] = MEM[1663] + MEM[2782];
assign MEM[15636] = MEM[1669] + MEM[5060];
assign MEM[15637] = MEM[1699] + MEM[10685];
assign MEM[15638] = MEM[1700] + MEM[9308];
assign MEM[15639] = MEM[1701] + MEM[10007];
assign MEM[15640] = MEM[1702] + MEM[15219];
assign MEM[15641] = MEM[1706] + MEM[11336];
assign MEM[15642] = MEM[1714] + MEM[1882];
assign MEM[15643] = MEM[1724] + MEM[9796];
assign MEM[15644] = MEM[1726] + MEM[11258];
assign MEM[15645] = MEM[1735] + MEM[11847];
assign MEM[15646] = MEM[1741] + MEM[8817];
assign MEM[15647] = MEM[1754] + MEM[10823];
assign MEM[15648] = MEM[1755] + MEM[9735];
assign MEM[15649] = MEM[1765] + MEM[11266];
assign MEM[15650] = MEM[1774] + MEM[9173];
assign MEM[15651] = MEM[1783] + MEM[9711];
assign MEM[15652] = MEM[1787] + MEM[9868];
assign MEM[15653] = MEM[1789] + MEM[13588];
assign MEM[15654] = MEM[1811] + MEM[3668];
assign MEM[15655] = MEM[1831] + MEM[12787];
assign MEM[15656] = MEM[1836] + MEM[4039];
assign MEM[15657] = MEM[1837] + MEM[11924];
assign MEM[15658] = MEM[1839] + MEM[11293];
assign MEM[15659] = MEM[1847] + MEM[13328];
assign MEM[15660] = MEM[1863] + MEM[5364];
assign MEM[15661] = MEM[1870] + MEM[9671];
assign MEM[15662] = MEM[1871] + MEM[9406];
assign MEM[15663] = MEM[1874] + MEM[11482];
assign MEM[15664] = MEM[1890] + MEM[7376];
assign MEM[15665] = MEM[1894] + MEM[11225];
assign MEM[15666] = MEM[1906] + MEM[10314];
assign MEM[15667] = MEM[1911] + MEM[13630];
assign MEM[15668] = MEM[1916] + MEM[11733];
assign MEM[15669] = MEM[1919] + MEM[10319];
assign MEM[15670] = MEM[1926] + MEM[12754];
assign MEM[15671] = MEM[1941] + MEM[1853];
assign MEM[15672] = MEM[1941] + MEM[9499];
assign MEM[15673] = MEM[1959] + MEM[9156];
assign MEM[15674] = MEM[1963] + MEM[9201];
assign MEM[15675] = MEM[1973] + MEM[11312];
assign MEM[15676] = MEM[1974] + MEM[8166];
assign MEM[15677] = MEM[1987] + MEM[9403];
assign MEM[15678] = MEM[1996] + MEM[11335];
assign MEM[15679] = MEM[2012] + MEM[9476];
assign MEM[15680] = MEM[2027] + MEM[10638];
assign MEM[15681] = MEM[2028] + MEM[11610];
assign MEM[15682] = MEM[2030] + MEM[8924];
assign MEM[15683] = MEM[2044] + MEM[10482];
assign MEM[15684] = MEM[2055] + MEM[11281];
assign MEM[15685] = MEM[2061] + MEM[7308];
assign MEM[15686] = MEM[2063] + MEM[7961];
assign MEM[15687] = MEM[2069] + MEM[9649];
assign MEM[15688] = MEM[2079] + MEM[9669];
assign MEM[15689] = MEM[2085] + MEM[8771];
assign MEM[15690] = MEM[2103] + MEM[7503];
assign MEM[15691] = MEM[2110] + MEM[10103];
assign MEM[15692] = MEM[2119] + MEM[14896];
assign MEM[15693] = MEM[2122] + MEM[2146];
assign MEM[15694] = MEM[2132] + MEM[10204];
assign MEM[15695] = MEM[2143] + MEM[12868];
assign MEM[15696] = MEM[2149] + MEM[9535];
assign MEM[15697] = MEM[2151] + MEM[11755];
assign MEM[15698] = MEM[2154] + MEM[11687];
assign MEM[15699] = MEM[2155] + MEM[9046];
assign MEM[15700] = MEM[2156] + MEM[6592];
assign MEM[15701] = MEM[2162] + MEM[9599];
assign MEM[15702] = MEM[2166] + MEM[12806];
assign MEM[15703] = MEM[2174] + MEM[11839];
assign MEM[15704] = MEM[2187] + MEM[3242];
assign MEM[15705] = MEM[2189] + MEM[10086];
assign MEM[15706] = MEM[2190] + MEM[9619];
assign MEM[15707] = MEM[2196] + MEM[10582];
assign MEM[15708] = MEM[2197] + MEM[2164];
assign MEM[15709] = MEM[2202] + MEM[15380];
assign MEM[15710] = MEM[2205] + MEM[12359];
assign MEM[15711] = MEM[2218] + MEM[11811];
assign MEM[15712] = MEM[2219] + MEM[11573];
assign MEM[15713] = MEM[2253] + MEM[11712];
assign MEM[15714] = MEM[2254] + MEM[12954];
assign MEM[15715] = MEM[2259] + MEM[11529];
assign MEM[15716] = MEM[2262] + MEM[9080];
assign MEM[15717] = MEM[2263] + MEM[10721];
assign MEM[15718] = MEM[2266] + MEM[6363];
assign MEM[15719] = MEM[2283] + MEM[11402];
assign MEM[15720] = MEM[2284] + MEM[13531];
assign MEM[15721] = MEM[2290] + MEM[4445];
assign MEM[15722] = MEM[2300] + MEM[11274];
assign MEM[15723] = MEM[2306] + MEM[11937];
assign MEM[15724] = MEM[2325] + MEM[8568];
assign MEM[15725] = MEM[2333] + MEM[9986];
assign MEM[15726] = MEM[2339] + MEM[10491];
assign MEM[15727] = MEM[2340] + MEM[13849];
assign MEM[15728] = MEM[2346] + MEM[11093];
assign MEM[15729] = MEM[2363] + MEM[7112];
assign MEM[15730] = MEM[2366] + MEM[9166];
assign MEM[15731] = MEM[2390] + MEM[11386];
assign MEM[15732] = MEM[2399] + MEM[10479];
assign MEM[15733] = MEM[2406] + MEM[9504];
assign MEM[15734] = MEM[2407] + MEM[6324];
assign MEM[15735] = MEM[2412] + MEM[5926];
assign MEM[15736] = MEM[2414] + MEM[11223];
assign MEM[15737] = MEM[2423] + MEM[11359];
assign MEM[15738] = MEM[2436] + MEM[3341];
assign MEM[15739] = MEM[2439] + MEM[11308];
assign MEM[15740] = MEM[2455] + MEM[12120];
assign MEM[15741] = MEM[2461] + MEM[8700];
assign MEM[15742] = MEM[2476] + MEM[8715];
assign MEM[15743] = MEM[2484] + MEM[11485];
assign MEM[15744] = MEM[2486] + MEM[6615];
assign MEM[15745] = MEM[2490] + MEM[8774];
assign MEM[15746] = MEM[2492] + MEM[15385];
assign MEM[15747] = MEM[2498] + MEM[9817];
assign MEM[15748] = MEM[2501] + MEM[3203];
assign MEM[15749] = MEM[2503] + MEM[10092];
assign MEM[15750] = MEM[2515] + MEM[3181];
assign MEM[15751] = MEM[2515] + MEM[12483];
assign MEM[15752] = MEM[2518] + MEM[11351];
assign MEM[15753] = MEM[2522] + MEM[7117];
assign MEM[15754] = MEM[2535] + MEM[11186];
assign MEM[15755] = MEM[2549] + MEM[7765];
assign MEM[15756] = MEM[2551] + MEM[11273];
assign MEM[15757] = MEM[2572] + MEM[11986];
assign MEM[15758] = MEM[2575] + MEM[10462];
assign MEM[15759] = MEM[2579] + MEM[8308];
assign MEM[15760] = MEM[2580] + MEM[12998];
assign MEM[15761] = MEM[2590] + MEM[10030];
assign MEM[15762] = MEM[2597] + MEM[2672];
assign MEM[15763] = MEM[2602] + MEM[6742];
assign MEM[15764] = MEM[2603] + MEM[11392];
assign MEM[15765] = MEM[2619] + MEM[8492];
assign MEM[15766] = MEM[2621] + MEM[12056];
assign MEM[15767] = MEM[2626] + MEM[2708];
assign MEM[15768] = MEM[2629] + MEM[9844];
assign MEM[15769] = MEM[2634] + MEM[11915];
assign MEM[15770] = MEM[2654] + MEM[9840];
assign MEM[15771] = MEM[2664] + MEM[11677];
assign MEM[15772] = MEM[2665] + MEM[5952];
assign MEM[15773] = MEM[2695] + MEM[3071];
assign MEM[15774] = MEM[2707] + MEM[7849];
assign MEM[15775] = MEM[2709] + MEM[2983];
assign MEM[15776] = MEM[2719] + MEM[14930];
assign MEM[15777] = MEM[2725] + MEM[9360];
assign MEM[15778] = MEM[2731] + MEM[15351];
assign MEM[15779] = MEM[2732] + MEM[10226];
assign MEM[15780] = MEM[2733] + MEM[6663];
assign MEM[15781] = MEM[2743] + MEM[11920];
assign MEM[15782] = MEM[2763] + MEM[8171];
assign MEM[15783] = MEM[2771] + MEM[9667];
assign MEM[15784] = MEM[2773] + MEM[10470];
assign MEM[15785] = MEM[2775] + MEM[7462];
assign MEM[15786] = MEM[2780] + MEM[9866];
assign MEM[15787] = MEM[2804] + MEM[5821];
assign MEM[15788] = MEM[2826] + MEM[11842];
assign MEM[15789] = MEM[2830] + MEM[10952];
assign MEM[15790] = MEM[2835] + MEM[10372];
assign MEM[15791] = MEM[2846] + MEM[9449];
assign MEM[15792] = MEM[2847] + MEM[5589];
assign MEM[15793] = MEM[2852] + MEM[9438];
assign MEM[15794] = MEM[2858] + MEM[9177];
assign MEM[15795] = MEM[2863] + MEM[10556];
assign MEM[15796] = MEM[2879] + MEM[11763];
assign MEM[15797] = MEM[2884] + MEM[6409];
assign MEM[15798] = MEM[2895] + MEM[8800];
assign MEM[15799] = MEM[2903] + MEM[11412];
assign MEM[15800] = MEM[2909] + MEM[11174];
assign MEM[15801] = MEM[2910] + MEM[11559];
assign MEM[15802] = MEM[2939] + MEM[9571];
assign MEM[15803] = MEM[2951] + MEM[9872];
assign MEM[15804] = MEM[2954] + MEM[12279];
assign MEM[15805] = MEM[2956] + MEM[8944];
assign MEM[15806] = MEM[2958] + MEM[10580];
assign MEM[15807] = MEM[2964] + MEM[8841];
assign MEM[15808] = MEM[2978] + MEM[4846];
assign MEM[15809] = MEM[2978] + MEM[11388];
assign MEM[15810] = MEM[2980] + MEM[3322];
assign MEM[15811] = MEM[2982] + MEM[10169];
assign MEM[15812] = MEM[2990] + MEM[11756];
assign MEM[15813] = MEM[2991] + MEM[10506];
assign MEM[15814] = MEM[3005] + MEM[10174];
assign MEM[15815] = MEM[3010] + MEM[13813];
assign MEM[15816] = MEM[3013] + MEM[6820];
assign MEM[15817] = MEM[3030] + MEM[9106];
assign MEM[15818] = MEM[3037] + MEM[10178];
assign MEM[15819] = MEM[3045] + MEM[10298];
assign MEM[15820] = MEM[3058] + MEM[14147];
assign MEM[15821] = MEM[3070] + MEM[13577];
assign MEM[15822] = MEM[3077] + MEM[142];
assign MEM[15823] = MEM[3079] + MEM[9852];
assign MEM[15824] = MEM[3087] + MEM[9015];
assign MEM[15825] = MEM[3098] + MEM[7904];
assign MEM[15826] = MEM[3106] + MEM[11138];
assign MEM[15827] = MEM[3117] + MEM[11300];
assign MEM[15828] = MEM[3131] + MEM[11328];
assign MEM[15829] = MEM[3135] + MEM[10048];
assign MEM[15830] = MEM[3142] + MEM[6567];
assign MEM[15831] = MEM[3172] + MEM[13818];
assign MEM[15832] = MEM[3173] + MEM[9643];
assign MEM[15833] = MEM[3183] + MEM[10396];
assign MEM[15834] = MEM[3194] + MEM[8136];
assign MEM[15835] = MEM[3194] + MEM[11121];
assign MEM[15836] = MEM[3198] + MEM[11216];
assign MEM[15837] = MEM[3228] + MEM[11974];
assign MEM[15838] = MEM[3234] + MEM[10523];
assign MEM[15839] = MEM[3263] + MEM[14501];
assign MEM[15840] = MEM[3266] + MEM[9564];
assign MEM[15841] = MEM[3293] + MEM[11196];
assign MEM[15842] = MEM[3294] + MEM[10089];
assign MEM[15843] = MEM[3299] + MEM[3814];
assign MEM[15844] = MEM[3315] + MEM[9455];
assign MEM[15845] = MEM[3318] + MEM[4234];
assign MEM[15846] = MEM[3325] + MEM[9415];
assign MEM[15847] = MEM[3335] + MEM[10603];
assign MEM[15848] = MEM[3343] + MEM[11891];
assign MEM[15849] = MEM[3348] + MEM[8213];
assign MEM[15850] = MEM[3351] + MEM[8026];
assign MEM[15851] = MEM[3375] + MEM[10682];
assign MEM[15852] = MEM[3379] + MEM[4263];
assign MEM[15853] = MEM[3381] + MEM[10211];
assign MEM[15854] = MEM[3386] + MEM[9875];
assign MEM[15855] = MEM[3388] + MEM[11197];
assign MEM[15856] = MEM[3390] + MEM[11181];
assign MEM[15857] = MEM[3398] + MEM[11025];
assign MEM[15858] = MEM[3407] + MEM[7566];
assign MEM[15859] = MEM[3411] + MEM[10869];
assign MEM[15860] = MEM[3418] + MEM[7337];
assign MEM[15861] = MEM[3419] + MEM[12981];
assign MEM[15862] = MEM[3426] + MEM[11343];
assign MEM[15863] = MEM[3428] + MEM[6269];
assign MEM[15864] = MEM[3430] + MEM[12467];
assign MEM[15865] = MEM[3436] + MEM[7917];
assign MEM[15866] = MEM[3455] + MEM[12158];
assign MEM[15867] = MEM[3462] + MEM[14013];
assign MEM[15868] = MEM[3468] + MEM[11876];
assign MEM[15869] = MEM[3471] + MEM[3891];
assign MEM[15870] = MEM[3482] + MEM[5290];
assign MEM[15871] = MEM[3491] + MEM[14873];
assign MEM[15872] = MEM[3492] + MEM[14871];
assign MEM[15873] = MEM[3524] + MEM[11522];
assign MEM[15874] = MEM[3527] + MEM[11084];
assign MEM[15875] = MEM[3534] + MEM[5206];
assign MEM[15876] = MEM[3541] + MEM[11927];
assign MEM[15877] = MEM[3558] + MEM[4847];
assign MEM[15878] = MEM[3559] + MEM[9273];
assign MEM[15879] = MEM[3589] + MEM[10166];
assign MEM[15880] = MEM[3590] + MEM[8998];
assign MEM[15881] = MEM[3603] + MEM[5710];
assign MEM[15882] = MEM[3615] + MEM[4194];
assign MEM[15883] = MEM[3631] + MEM[9928];
assign MEM[15884] = MEM[3635] + MEM[8866];
assign MEM[15885] = MEM[3644] + MEM[7574];
assign MEM[15886] = MEM[3650] + MEM[10138];
assign MEM[15887] = MEM[3651] + MEM[10739];
assign MEM[15888] = MEM[3662] + MEM[7320];
assign MEM[15889] = MEM[3692] + MEM[12575];
assign MEM[15890] = MEM[3693] + MEM[8745];
assign MEM[15891] = MEM[3699] + MEM[12403];
assign MEM[15892] = MEM[3700] + MEM[10112];
assign MEM[15893] = MEM[3701] + MEM[8798];
assign MEM[15894] = MEM[3749] + MEM[13224];
assign MEM[15895] = MEM[3751] + MEM[13490];
assign MEM[15896] = MEM[3765] + MEM[11521];
assign MEM[15897] = MEM[3791] + MEM[7017];
assign MEM[15898] = MEM[3821] + MEM[11567];
assign MEM[15899] = MEM[3826] + MEM[5814];
assign MEM[15900] = MEM[3838] + MEM[8876];
assign MEM[15901] = MEM[3843] + MEM[10619];
assign MEM[15902] = MEM[3844] + MEM[11425];
assign MEM[15903] = MEM[3851] + MEM[12655];
assign MEM[15904] = MEM[3852] + MEM[7478];
assign MEM[15905] = MEM[3862] + MEM[13427];
assign MEM[15906] = MEM[3875] + MEM[10006];
assign MEM[15907] = MEM[3878] + MEM[12880];
assign MEM[15908] = MEM[3882] + MEM[6499];
assign MEM[15909] = MEM[3894] + MEM[11597];
assign MEM[15910] = MEM[3917] + MEM[9297];
assign MEM[15911] = MEM[3919] + MEM[11280];
assign MEM[15912] = MEM[3922] + MEM[10375];
assign MEM[15913] = MEM[3927] + MEM[9950];
assign MEM[15914] = MEM[3932] + MEM[4061];
assign MEM[15915] = MEM[3934] + MEM[11342];
assign MEM[15916] = MEM[3935] + MEM[11476];
assign MEM[15917] = MEM[3954] + MEM[9988];
assign MEM[15918] = MEM[3966] + MEM[9971];
assign MEM[15919] = MEM[3982] + MEM[9167];
assign MEM[15920] = MEM[3986] + MEM[8988];
assign MEM[15921] = MEM[3990] + MEM[11510];
assign MEM[15922] = MEM[3991] + MEM[9674];
assign MEM[15923] = MEM[4029] + MEM[2790];
assign MEM[15924] = MEM[4055] + MEM[11908];
assign MEM[15925] = MEM[4061] + MEM[12845];
assign MEM[15926] = MEM[4063] + MEM[10825];
assign MEM[15927] = MEM[4068] + MEM[11291];
assign MEM[15928] = MEM[4071] + MEM[12789];
assign MEM[15929] = MEM[4084] + MEM[5701];
assign MEM[15930] = MEM[4101] + MEM[6798];
assign MEM[15931] = MEM[4114] + MEM[13990];
assign MEM[15932] = MEM[4125] + MEM[11747];
assign MEM[15933] = MEM[4139] + MEM[9547];
assign MEM[15934] = MEM[4149] + MEM[9725];
assign MEM[15935] = MEM[4173] + MEM[11390];
assign MEM[15936] = MEM[4181] + MEM[13537];
assign MEM[15937] = MEM[4204] + MEM[11133];
assign MEM[15938] = MEM[4205] + MEM[11292];
assign MEM[15939] = MEM[4213] + MEM[6369];
assign MEM[15940] = MEM[4215] + MEM[8393];
assign MEM[15941] = MEM[4220] + MEM[11745];
assign MEM[15942] = MEM[4226] + MEM[5947];
assign MEM[15943] = MEM[4239] + MEM[7208];
assign MEM[15944] = MEM[4247] + MEM[9791];
assign MEM[15945] = MEM[4251] + MEM[10483];
assign MEM[15946] = MEM[4253] + MEM[11593];
assign MEM[15947] = MEM[4255] + MEM[10188];
assign MEM[15948] = MEM[4269] + MEM[14868];
assign MEM[15949] = MEM[4275] + MEM[8207];
assign MEM[15950] = MEM[4277] + MEM[4634];
assign MEM[15951] = MEM[4279] + MEM[11398];
assign MEM[15952] = MEM[4295] + MEM[11233];
assign MEM[15953] = MEM[4301] + MEM[9313];
assign MEM[15954] = MEM[4303] + MEM[10097];
assign MEM[15955] = MEM[4317] + MEM[5459];
assign MEM[15956] = MEM[4330] + MEM[2999];
assign MEM[15957] = MEM[4331] + MEM[9320];
assign MEM[15958] = MEM[4348] + MEM[8394];
assign MEM[15959] = MEM[4362] + MEM[5381];
assign MEM[15960] = MEM[4364] + MEM[12178];
assign MEM[15961] = MEM[4365] + MEM[12275];
assign MEM[15962] = MEM[4383] + MEM[11841];
assign MEM[15963] = MEM[4391] + MEM[8028];
assign MEM[15964] = MEM[4395] + MEM[9931];
assign MEM[15965] = MEM[4397] + MEM[9365];
assign MEM[15966] = MEM[4402] + MEM[5110];
assign MEM[15967] = MEM[4403] + MEM[10170];
assign MEM[15968] = MEM[4404] + MEM[11987];
assign MEM[15969] = MEM[4411] + MEM[11093];
assign MEM[15970] = MEM[4434] + MEM[8245];
assign MEM[15971] = MEM[4444] + MEM[7995];
assign MEM[15972] = MEM[4458] + MEM[10275];
assign MEM[15973] = MEM[4485] + MEM[11220];
assign MEM[15974] = MEM[4498] + MEM[12653];
assign MEM[15975] = MEM[4510] + MEM[11249];
assign MEM[15976] = MEM[4516] + MEM[10132];
assign MEM[15977] = MEM[4527] + MEM[10490];
assign MEM[15978] = MEM[4533] + MEM[11535];
assign MEM[15979] = MEM[4534] + MEM[10445];
assign MEM[15980] = MEM[4549] + MEM[9584];
assign MEM[15981] = MEM[4550] + MEM[11132];
assign MEM[15982] = MEM[4558] + MEM[10385];
assign MEM[15983] = MEM[4566] + MEM[11527];
assign MEM[15984] = MEM[4571] + MEM[13740];
assign MEM[15985] = MEM[4574] + MEM[11102];
assign MEM[15986] = MEM[4575] + MEM[11302];
assign MEM[15987] = MEM[4596] + MEM[11822];
assign MEM[15988] = MEM[4597] + MEM[11345];
assign MEM[15989] = MEM[4610] + MEM[15301];
assign MEM[15990] = MEM[4635] + MEM[9092];
assign MEM[15991] = MEM[4636] + MEM[11506];
assign MEM[15992] = MEM[4638] + MEM[11461];
assign MEM[15993] = MEM[4646] + MEM[9175];
assign MEM[15994] = MEM[4650] + MEM[15361];
assign MEM[15995] = MEM[4666] + MEM[9589];
assign MEM[15996] = MEM[4668] + MEM[11387];
assign MEM[15997] = MEM[4670] + MEM[11451];
assign MEM[15998] = MEM[4682] + MEM[12830];
assign MEM[15999] = MEM[4733] + MEM[11519];
assign MEM[16000] = MEM[4735] + MEM[5486];
assign MEM[16001] = MEM[4740] + MEM[11404];
assign MEM[16002] = MEM[4743] + MEM[5682];
assign MEM[16003] = MEM[4758] + MEM[12112];
assign MEM[16004] = MEM[4763] + MEM[11836];
assign MEM[16005] = MEM[4771] + MEM[10866];
assign MEM[16006] = MEM[4773] + MEM[7622];
assign MEM[16007] = MEM[4794] + MEM[14772];
assign MEM[16008] = MEM[4813] + MEM[11759];
assign MEM[16009] = MEM[4831] + MEM[9908];
assign MEM[16010] = MEM[4859] + MEM[11362];
assign MEM[16011] = MEM[4860] + MEM[4591];
assign MEM[16012] = MEM[4866] + MEM[13369];
assign MEM[16013] = MEM[4874] + MEM[10737];
assign MEM[16014] = MEM[4892] + MEM[11418];
assign MEM[16015] = MEM[4894] + MEM[10318];
assign MEM[16016] = MEM[4902] + MEM[9883];
assign MEM[16017] = MEM[4906] + MEM[8078];
assign MEM[16018] = MEM[4918] + MEM[10227];
assign MEM[16019] = MEM[4946] + MEM[9514];
assign MEM[16020] = MEM[4956] + MEM[11232];
assign MEM[16021] = MEM[4963] + MEM[10104];
assign MEM[16022] = MEM[4973] + MEM[9737];
assign MEM[16023] = MEM[4979] + MEM[8083];
assign MEM[16024] = MEM[4997] + MEM[7123];
assign MEM[16025] = MEM[5015] + MEM[9733];
assign MEM[16026] = MEM[5027] + MEM[12960];
assign MEM[16027] = MEM[5029] + MEM[10144];
assign MEM[16028] = MEM[5037] + MEM[7098];
assign MEM[16029] = MEM[5039] + MEM[8967];
assign MEM[16030] = MEM[5050] + MEM[11534];
assign MEM[16031] = MEM[5062] + MEM[9500];
assign MEM[16032] = MEM[5077] + MEM[11311];
assign MEM[16033] = MEM[5082] + MEM[9059];
assign MEM[16034] = MEM[5092] + MEM[11465];
assign MEM[16035] = MEM[5101] + MEM[13768];
assign MEM[16036] = MEM[5107] + MEM[11523];
assign MEM[16037] = MEM[5114] + MEM[10745];
assign MEM[16038] = MEM[5118] + MEM[9542];
assign MEM[16039] = MEM[5134] + MEM[10025];
assign MEM[16040] = MEM[5141] + MEM[10016];
assign MEM[16041] = MEM[5158] + MEM[12827];
assign MEM[16042] = MEM[5159] + MEM[8976];
assign MEM[16043] = MEM[5165] + MEM[8462];
assign MEM[16044] = MEM[5166] + MEM[10790];
assign MEM[16045] = MEM[5179] + MEM[11151];
assign MEM[16046] = MEM[5182] + MEM[10980];
assign MEM[16047] = MEM[5189] + MEM[11898];
assign MEM[16048] = MEM[5190] + MEM[9215];
assign MEM[16049] = MEM[5194] + MEM[9316];
assign MEM[16050] = MEM[5212] + MEM[6023];
assign MEM[16051] = MEM[5215] + MEM[12914];
assign MEM[16052] = MEM[5231] + MEM[4604];
assign MEM[16053] = MEM[5238] + MEM[11505];
assign MEM[16054] = MEM[5244] + MEM[10545];
assign MEM[16055] = MEM[5262] + MEM[13338];
assign MEM[16056] = MEM[5275] + MEM[9717];
assign MEM[16057] = MEM[5309] + MEM[12111];
assign MEM[16058] = MEM[5312] + MEM[9544];
assign MEM[16059] = MEM[5323] + MEM[13122];
assign MEM[16060] = MEM[5325] + MEM[6376];
assign MEM[16061] = MEM[5332] + MEM[10489];
assign MEM[16062] = MEM[5340] + MEM[7034];
assign MEM[16063] = MEM[5341] + MEM[11373];
assign MEM[16064] = MEM[5358] + MEM[8132];
assign MEM[16065] = MEM[5359] + MEM[9565];
assign MEM[16066] = MEM[5375] + MEM[9646];
assign MEM[16067] = MEM[5390] + MEM[12724];
assign MEM[16068] = MEM[5391] + MEM[11949];
assign MEM[16069] = MEM[5397] + MEM[6545];
assign MEM[16070] = MEM[5410] + MEM[9263];
assign MEM[16071] = MEM[5415] + MEM[11349];
assign MEM[16072] = MEM[5422] + MEM[11829];
assign MEM[16073] = MEM[5423] + MEM[10863];
assign MEM[16074] = MEM[5431] + MEM[8337];
assign MEM[16075] = MEM[5436] + MEM[9886];
assign MEM[16076] = MEM[5453] + MEM[11511];
assign MEM[16077] = MEM[5454] + MEM[8918];
assign MEM[16078] = MEM[5455] + MEM[11565];
assign MEM[16079] = MEM[5460] + MEM[7284];
assign MEM[16080] = MEM[5484] + MEM[9946];
assign MEM[16081] = MEM[5485] + MEM[11095];
assign MEM[16082] = MEM[5491] + MEM[7356];
assign MEM[16083] = MEM[5494] + MEM[6196];
assign MEM[16084] = MEM[5502] + MEM[9724];
assign MEM[16085] = MEM[5511] + MEM[8235];
assign MEM[16086] = MEM[5514] + MEM[10393];
assign MEM[16087] = MEM[5517] + MEM[10126];
assign MEM[16088] = MEM[5535] + MEM[6897];
assign MEM[16089] = MEM[5538] + MEM[9707];
assign MEM[16090] = MEM[5543] + MEM[9841];
assign MEM[16091] = MEM[5547] + MEM[11655];
assign MEM[16092] = MEM[5550] + MEM[10214];
assign MEM[16093] = MEM[5554] + MEM[11922];
assign MEM[16094] = MEM[5556] + MEM[10201];
assign MEM[16095] = MEM[5565] + MEM[7872];
assign MEM[16096] = MEM[5597] + MEM[10801];
assign MEM[16097] = MEM[5599] + MEM[10315];
assign MEM[16098] = MEM[5607] + MEM[10573];
assign MEM[16099] = MEM[5613] + MEM[10133];
assign MEM[16100] = MEM[5631] + MEM[15190];
assign MEM[16101] = MEM[5660] + MEM[9755];
assign MEM[16102] = MEM[5667] + MEM[11997];
assign MEM[16103] = MEM[5669] + MEM[3372];
assign MEM[16104] = MEM[5685] + MEM[12890];
assign MEM[16105] = MEM[5687] + MEM[9703];
assign MEM[16106] = MEM[5691] + MEM[10636];
assign MEM[16107] = MEM[5707] + MEM[10291];
assign MEM[16108] = MEM[5714] + MEM[7843];
assign MEM[16109] = MEM[5716] + MEM[14559];
assign MEM[16110] = MEM[5719] + MEM[12255];
assign MEM[16111] = MEM[5734] + MEM[12641];
assign MEM[16112] = MEM[5739] + MEM[11301];
assign MEM[16113] = MEM[5758] + MEM[12190];
assign MEM[16114] = MEM[5764] + MEM[11467];
assign MEM[16115] = MEM[5775] + MEM[8224];
assign MEM[16116] = MEM[5795] + MEM[6784];
assign MEM[16117] = MEM[5796] + MEM[9862];
assign MEM[16118] = MEM[5831] + MEM[12687];
assign MEM[16119] = MEM[5853] + MEM[11151];
assign MEM[16120] = MEM[5877] + MEM[6446];
assign MEM[16121] = MEM[5887] + MEM[11415];
assign MEM[16122] = MEM[5893] + MEM[10295];
assign MEM[16123] = MEM[5898] + MEM[11318];
assign MEM[16124] = MEM[5907] + MEM[11769];
assign MEM[16125] = MEM[5915] + MEM[9926];
assign MEM[16126] = MEM[5916] + MEM[9600];
assign MEM[16127] = MEM[5917] + MEM[12094];
assign MEM[16128] = MEM[5918] + MEM[11278];
assign MEM[16129] = MEM[5950] + MEM[11326];
assign MEM[16130] = MEM[5951] + MEM[10184];
assign MEM[16131] = MEM[5953] + MEM[11856];
assign MEM[16132] = MEM[5957] + MEM[6902];
assign MEM[16133] = MEM[5958] + MEM[11352];
assign MEM[16134] = MEM[5966] + MEM[11463];
assign MEM[16135] = MEM[6003] + MEM[11789];
assign MEM[16136] = MEM[6029] + MEM[13251];
assign MEM[16137] = MEM[6061] + MEM[5444];
assign MEM[16138] = MEM[6086] + MEM[10583];
assign MEM[16139] = MEM[6101] + MEM[10255];
assign MEM[16140] = MEM[6108] + MEM[9540];
assign MEM[16141] = MEM[6118] + MEM[9774];
assign MEM[16142] = MEM[6131] + MEM[12434];
assign MEM[16143] = MEM[6150] + MEM[12547];
assign MEM[16144] = MEM[6164] + MEM[10244];
assign MEM[16145] = MEM[6166] + MEM[9884];
assign MEM[16146] = MEM[6188] + MEM[10284];
assign MEM[16147] = MEM[6189] + MEM[12661];
assign MEM[16148] = MEM[6197] + MEM[11344];
assign MEM[16149] = MEM[6212] + MEM[7280];
assign MEM[16150] = MEM[6239] + MEM[9022];
assign MEM[16151] = MEM[6246] + MEM[7184];
assign MEM[16152] = MEM[6247] + MEM[11460];
assign MEM[16153] = MEM[6271] + MEM[12338];
assign MEM[16154] = MEM[6272] + MEM[9104];
assign MEM[16155] = MEM[6288] + MEM[11694];
assign MEM[16156] = MEM[6296] + MEM[11221];
assign MEM[16157] = MEM[6304] + MEM[7496];
assign MEM[16158] = MEM[6305] + MEM[9640];
assign MEM[16159] = MEM[6318] + MEM[10026];
assign MEM[16160] = MEM[6330] + MEM[10587];
assign MEM[16161] = MEM[6334] + MEM[11179];
assign MEM[16162] = MEM[6341] + MEM[10137];
assign MEM[16163] = MEM[6342] + MEM[9783];
assign MEM[16164] = MEM[6359] + MEM[10236];
assign MEM[16165] = MEM[6361] + MEM[7178];
assign MEM[16166] = MEM[6373] + MEM[6843];
assign MEM[16167] = MEM[6374] + MEM[11854];
assign MEM[16168] = MEM[6381] + MEM[10564];
assign MEM[16169] = MEM[6388] + MEM[11309];
assign MEM[16170] = MEM[6405] + MEM[12266];
assign MEM[16171] = MEM[6411] + MEM[10610];
assign MEM[16172] = MEM[6413] + MEM[11555];
assign MEM[16173] = MEM[6453] + MEM[10536];
assign MEM[16174] = MEM[6470] + MEM[6977];
assign MEM[16175] = MEM[6494] + MEM[9574];
assign MEM[16176] = MEM[6514] + MEM[11085];
assign MEM[16177] = MEM[6515] + MEM[8049];
assign MEM[16178] = MEM[6516] + MEM[9801];
assign MEM[16179] = MEM[6518] + MEM[12055];
assign MEM[16180] = MEM[6532] + MEM[10539];
assign MEM[16181] = MEM[6534] + MEM[10142];
assign MEM[16182] = MEM[6537] + MEM[7312];
assign MEM[16183] = MEM[6557] + MEM[12952];
assign MEM[16184] = MEM[6558] + MEM[7128];
assign MEM[16185] = MEM[6569] + MEM[9821];
assign MEM[16186] = MEM[6578] + MEM[11985];
assign MEM[16187] = MEM[6585] + MEM[11831];
assign MEM[16188] = MEM[6592] + MEM[13802];
assign MEM[16189] = MEM[6597] + MEM[11426];
assign MEM[16190] = MEM[6606] + MEM[6906];
assign MEM[16191] = MEM[6610] + MEM[11456];
assign MEM[16192] = MEM[6614] + MEM[7532];
assign MEM[16193] = MEM[6619] + MEM[10113];
assign MEM[16194] = MEM[6651] + MEM[9009];
assign MEM[16195] = MEM[6662] + MEM[13234];
assign MEM[16196] = MEM[6677] + MEM[8741];
assign MEM[16197] = MEM[6737] + MEM[7255];
assign MEM[16198] = MEM[6739] + MEM[6879];
assign MEM[16199] = MEM[6746] + MEM[9481];
assign MEM[16200] = MEM[6755] + MEM[9876];
assign MEM[16201] = MEM[6779] + MEM[9705];
assign MEM[16202] = MEM[6800] + MEM[8503];
assign MEM[16203] = MEM[6801] + MEM[11340];
assign MEM[16204] = MEM[6806] + MEM[9361];
assign MEM[16205] = MEM[6807] + MEM[13124];
assign MEM[16206] = MEM[6808] + MEM[11533];
assign MEM[16207] = MEM[6818] + MEM[9681];
assign MEM[16208] = MEM[6822] + MEM[11256];
assign MEM[16209] = MEM[6839] + MEM[11428];
assign MEM[16210] = MEM[6855] + MEM[9803];
assign MEM[16211] = MEM[6856] + MEM[11667];
assign MEM[16212] = MEM[6857] + MEM[11823];
assign MEM[16213] = MEM[6876] + MEM[9314];
assign MEM[16214] = MEM[6885] + MEM[10377];
assign MEM[16215] = MEM[6893] + MEM[11940];
assign MEM[16216] = MEM[6898] + MEM[10744];
assign MEM[16217] = MEM[6909] + MEM[11724];
assign MEM[16218] = MEM[6911] + MEM[12866];
assign MEM[16219] = MEM[6912] + MEM[12978];
assign MEM[16220] = MEM[6913] + MEM[6022];
assign MEM[16221] = MEM[6917] + MEM[13458];
assign MEM[16222] = MEM[6930] + MEM[10259];
assign MEM[16223] = MEM[6937] + MEM[11598];
assign MEM[16224] = MEM[6945] + MEM[11853];
assign MEM[16225] = MEM[6960] + MEM[11089];
assign MEM[16226] = MEM[6966] + MEM[9936];
assign MEM[16227] = MEM[6980] + MEM[7035];
assign MEM[16228] = MEM[6986] + MEM[13462];
assign MEM[16229] = MEM[7004] + MEM[13352];
assign MEM[16230] = MEM[7024] + MEM[11276];
assign MEM[16231] = MEM[7027] + MEM[9804];
assign MEM[16232] = MEM[7030] + MEM[10513];
assign MEM[16233] = MEM[7033] + MEM[10543];
assign MEM[16234] = MEM[7036] + MEM[12193];
assign MEM[16235] = MEM[7047] + MEM[4645];
assign MEM[16236] = MEM[7049] + MEM[10562];
assign MEM[16237] = MEM[7057] + MEM[11843];
assign MEM[16238] = MEM[7059] + MEM[9330];
assign MEM[16239] = MEM[7074] + MEM[9392];
assign MEM[16240] = MEM[7075] + MEM[10069];
assign MEM[16241] = MEM[7095] + MEM[11433];
assign MEM[16242] = MEM[7104] + MEM[9090];
assign MEM[16243] = MEM[7108] + MEM[11950];
assign MEM[16244] = MEM[7111] + MEM[11872];
assign MEM[16245] = MEM[7122] + MEM[11406];
assign MEM[16246] = MEM[7127] + MEM[13728];
assign MEM[16247] = MEM[7138] + MEM[12066];
assign MEM[16248] = MEM[7145] + MEM[12163];
assign MEM[16249] = MEM[7148] + MEM[5750];
assign MEM[16250] = MEM[7149] + MEM[10727];
assign MEM[16251] = MEM[7177] + MEM[12607];
assign MEM[16252] = MEM[7191] + MEM[12503];
assign MEM[16253] = MEM[7198] + MEM[10075];
assign MEM[16254] = MEM[7202] + MEM[9850];
assign MEM[16255] = MEM[7211] + MEM[9332];
assign MEM[16256] = MEM[7215] + MEM[10531];
assign MEM[16257] = MEM[7243] + MEM[9782];
assign MEM[16258] = MEM[7250] + MEM[9569];
assign MEM[16259] = MEM[7281] + MEM[10938];
assign MEM[16260] = MEM[7282] + MEM[10180];
assign MEM[16261] = MEM[7288] + MEM[3971];
assign MEM[16262] = MEM[7289] + MEM[11913];
assign MEM[16263] = MEM[7291] + MEM[8191];
assign MEM[16264] = MEM[7292] + MEM[10693];
assign MEM[16265] = MEM[7297] + MEM[9546];
assign MEM[16266] = MEM[7307] + MEM[11764];
assign MEM[16267] = MEM[7314] + MEM[11284];
assign MEM[16268] = MEM[7318] + MEM[10357];
assign MEM[16269] = MEM[7322] + MEM[10179];
assign MEM[16270] = MEM[7323] + MEM[11255];
assign MEM[16271] = MEM[7328] + MEM[10652];
assign MEM[16272] = MEM[7344] + MEM[9775];
assign MEM[16273] = MEM[7349] + MEM[5338];
assign MEM[16274] = MEM[7353] + MEM[10908];
assign MEM[16275] = MEM[7354] + MEM[11229];
assign MEM[16276] = MEM[7370] + MEM[11560];
assign MEM[16277] = MEM[7383] + MEM[10123];
assign MEM[16278] = MEM[7385] + MEM[10419];
assign MEM[16279] = MEM[7390] + MEM[9435];
assign MEM[16280] = MEM[7409] + MEM[11244];
assign MEM[16281] = MEM[7410] + MEM[10717];
assign MEM[16282] = MEM[7433] + MEM[9558];
assign MEM[16283] = MEM[7436] + MEM[11187];
assign MEM[16284] = MEM[7461] + MEM[8834];
assign MEM[16285] = MEM[7471] + MEM[11941];
assign MEM[16286] = MEM[7476] + MEM[6709];
assign MEM[16287] = MEM[7479] + MEM[9035];
assign MEM[16288] = MEM[7499] + MEM[11568];
assign MEM[16289] = MEM[7500] + MEM[8980];
assign MEM[16290] = MEM[7501] + MEM[14771];
assign MEM[16291] = MEM[7505] + MEM[3893];
assign MEM[16292] = MEM[7510] + MEM[11294];
assign MEM[16293] = MEM[7534] + MEM[10758];
assign MEM[16294] = MEM[7540] + MEM[11569];
assign MEM[16295] = MEM[7541] + MEM[10496];
assign MEM[16296] = MEM[7580] + MEM[11650];
assign MEM[16297] = MEM[7589] + MEM[10111];
assign MEM[16298] = MEM[7612] + MEM[10181];
assign MEM[16299] = MEM[7626] + MEM[10401];
assign MEM[16300] = MEM[7629] + MEM[8645];
assign MEM[16301] = MEM[7630] + MEM[8407];
assign MEM[16302] = MEM[7632] + MEM[9256];
assign MEM[16303] = MEM[7645] + MEM[5175];
assign MEM[16304] = MEM[7662] + MEM[11431];
assign MEM[16305] = MEM[7670] + MEM[11862];
assign MEM[16306] = MEM[7673] + MEM[10072];
assign MEM[16307] = MEM[7677] + MEM[11753];
assign MEM[16308] = MEM[7709] + MEM[12988];
assign MEM[16309] = MEM[7713] + MEM[9767];
assign MEM[16310] = MEM[7720] + MEM[11170];
assign MEM[16311] = MEM[7733] + MEM[9199];
assign MEM[16312] = MEM[7748] + MEM[12224];
assign MEM[16313] = MEM[7758] + MEM[9487];
assign MEM[16314] = MEM[7763] + MEM[11608];
assign MEM[16315] = MEM[7764] + MEM[11462];
assign MEM[16316] = MEM[7769] + MEM[10698];
assign MEM[16317] = MEM[7791] + MEM[11314];
assign MEM[16318] = MEM[7796] + MEM[11780];
assign MEM[16319] = MEM[7799] + MEM[11499];
assign MEM[16320] = MEM[7801] + MEM[6390];
assign MEM[16321] = MEM[7802] + MEM[11215];
assign MEM[16322] = MEM[7803] + MEM[9969];
assign MEM[16323] = MEM[7804] + MEM[10526];
assign MEM[16324] = MEM[7806] + MEM[11590];
assign MEM[16325] = MEM[7809] + MEM[9193];
assign MEM[16326] = MEM[7813] + MEM[12411];
assign MEM[16327] = MEM[7818] + MEM[8548];
assign MEM[16328] = MEM[7820] + MEM[11758];
assign MEM[16329] = MEM[7870] + MEM[11374];
assign MEM[16330] = MEM[7875] + MEM[8957];
assign MEM[16331] = MEM[7879] + MEM[9551];
assign MEM[16332] = MEM[7885] + MEM[9987];
assign MEM[16333] = MEM[7892] + MEM[11488];
assign MEM[16334] = MEM[7899] + MEM[10276];
assign MEM[16335] = MEM[7915] + MEM[11697];
assign MEM[16336] = MEM[7931] + MEM[9467];
assign MEM[16337] = MEM[7941] + MEM[8866];
assign MEM[16338] = MEM[7946] + MEM[12005];
assign MEM[16339] = MEM[7952] + MEM[9384];
assign MEM[16340] = MEM[7959] + MEM[10585];
assign MEM[16341] = MEM[7961] + MEM[13386];
assign MEM[16342] = MEM[7962] + MEM[6838];
assign MEM[16343] = MEM[7970] + MEM[13329];
assign MEM[16344] = MEM[7975] + MEM[10307];
assign MEM[16345] = MEM[7976] + MEM[10575];
assign MEM[16346] = MEM[7985] + MEM[10064];
assign MEM[16347] = MEM[7989] + MEM[10554];
assign MEM[16348] = MEM[7997] + MEM[8696];
assign MEM[16349] = MEM[7999] + MEM[11486];
assign MEM[16350] = MEM[8010] + MEM[9734];
assign MEM[16351] = MEM[8017] + MEM[10024];
assign MEM[16352] = MEM[8027] + MEM[10498];
assign MEM[16353] = MEM[8030] + MEM[12859];
assign MEM[16354] = MEM[8032] + MEM[10432];
assign MEM[16355] = MEM[8036] + MEM[8045];
assign MEM[16356] = MEM[8048] + MEM[8994];
assign MEM[16357] = MEM[8051] + MEM[10306];
assign MEM[16358] = MEM[8066] + MEM[6015];
assign MEM[16359] = MEM[8067] + MEM[13120];
assign MEM[16360] = MEM[8084] + MEM[8676];
assign MEM[16361] = MEM[8085] + MEM[9223];
assign MEM[16362] = MEM[8091] + MEM[9922];
assign MEM[16363] = MEM[8102] + MEM[10467];
assign MEM[16364] = MEM[8104] + MEM[12793];
assign MEM[16365] = MEM[8112] + MEM[10469];
assign MEM[16366] = MEM[8116] + MEM[8378];
assign MEM[16367] = MEM[8116] + MEM[9299];
assign MEM[16368] = MEM[8134] + MEM[11424];
assign MEM[16369] = MEM[8138] + MEM[13049];
assign MEM[16370] = MEM[8161] + MEM[12372];
assign MEM[16371] = MEM[8188] + MEM[12053];
assign MEM[16372] = MEM[8208] + MEM[9460];
assign MEM[16373] = MEM[8218] + MEM[9833];
assign MEM[16374] = MEM[8230] + MEM[8401];
assign MEM[16375] = MEM[8237] + MEM[10705];
assign MEM[16376] = MEM[8240] + MEM[10515];
assign MEM[16377] = MEM[8241] + MEM[10623];
assign MEM[16378] = MEM[8243] + MEM[13235];
assign MEM[16379] = MEM[8263] + MEM[11520];
assign MEM[16380] = MEM[8265] + MEM[11353];
assign MEM[16381] = MEM[8278] + MEM[6465];
assign MEM[16382] = MEM[8282] + MEM[8368];
assign MEM[16383] = MEM[8283] + MEM[9525];
assign MEM[16384] = MEM[8288] + MEM[12943];
assign MEM[16385] = MEM[8289] + MEM[12326];
assign MEM[16386] = MEM[8299] + MEM[11277];
assign MEM[16387] = MEM[8304] + MEM[11615];
assign MEM[16388] = MEM[8309] + MEM[11072];
assign MEM[16389] = MEM[8316] + MEM[12654];
assign MEM[16390] = MEM[8326] + MEM[11791];
assign MEM[16391] = MEM[8335] + MEM[13297];
assign MEM[16392] = MEM[8367] + MEM[10252];
assign MEM[16393] = MEM[8369] + MEM[11703];
assign MEM[16394] = MEM[8371] + MEM[11757];
assign MEM[16395] = MEM[8380] + MEM[9831];
assign MEM[16396] = MEM[8392] + MEM[12519];
assign MEM[16397] = MEM[8397] + MEM[9871];
assign MEM[16398] = MEM[8405] + MEM[10135];
assign MEM[16399] = MEM[8412] + MEM[11984];
assign MEM[16400] = MEM[8430] + MEM[10992];
assign MEM[16401] = MEM[8438] + MEM[8947];
assign MEM[16402] = MEM[8448] + MEM[14231];
assign MEM[16403] = MEM[8452] + MEM[10102];
assign MEM[16404] = MEM[8472] + MEM[12552];
assign MEM[16405] = MEM[8474] + MEM[11770];
assign MEM[16406] = MEM[8482] + MEM[9636];
assign MEM[16407] = MEM[8484] + MEM[11183];
assign MEM[16408] = MEM[8489] + MEM[13554];
assign MEM[16409] = MEM[8493] + MEM[13324];
assign MEM[16410] = MEM[8518] + MEM[10605];
assign MEM[16411] = MEM[8522] + MEM[9714];
assign MEM[16412] = MEM[8525] + MEM[9834];
assign MEM[16413] = MEM[8527] + MEM[9802];
assign MEM[16414] = MEM[8528] + MEM[9663];
assign MEM[16415] = MEM[8534] + MEM[12046];
assign MEM[16416] = MEM[8549] + MEM[10157];
assign MEM[16417] = MEM[8552] + MEM[8939];
assign MEM[16418] = MEM[8557] + MEM[11713];
assign MEM[16419] = MEM[8570] + MEM[11385];
assign MEM[16420] = MEM[8589] + MEM[9641];
assign MEM[16421] = MEM[8590] + MEM[12186];
assign MEM[16422] = MEM[8616] + MEM[12328];
assign MEM[16423] = MEM[8622] + MEM[10050];
assign MEM[16424] = MEM[8631] + MEM[8924];
assign MEM[16425] = MEM[8639] + MEM[13283];
assign MEM[16426] = MEM[8642] + MEM[11446];
assign MEM[16427] = MEM[8651] + MEM[6455];
assign MEM[16428] = MEM[8656] + MEM[11711];
assign MEM[16429] = MEM[8657] + MEM[10505];
assign MEM[16430] = MEM[8659] + MEM[12958];
assign MEM[16431] = MEM[8660] + MEM[12946];
assign MEM[16432] = MEM[8664] + MEM[9698];
assign MEM[16433] = MEM[8668] + MEM[10994];
assign MEM[16434] = MEM[8673] + MEM[10020];
assign MEM[16435] = MEM[8679] + MEM[16060];
assign MEM[16436] = MEM[8695] + MEM[9917];
assign MEM[16437] = MEM[8705] + MEM[10817];
assign MEM[16438] = MEM[8728] + MEM[11609];
assign MEM[16439] = MEM[8733] + MEM[11163];
assign MEM[16440] = MEM[8734] + MEM[7225];
assign MEM[16441] = MEM[8751] + MEM[7137];
assign MEM[16442] = MEM[8755] + MEM[10099];
assign MEM[16443] = MEM[8785] + MEM[9691];
assign MEM[16444] = MEM[8807] + MEM[11582];
assign MEM[16445] = MEM[8832] + MEM[14217];
assign MEM[16446] = MEM[8850] + MEM[9020];
assign MEM[16447] = MEM[8856] + MEM[10561];
assign MEM[16448] = MEM[8873] + MEM[9257];
assign MEM[16449] = MEM[8885] + MEM[10783];
assign MEM[16450] = MEM[8888] + MEM[10468];
assign MEM[16451] = MEM[8896] + MEM[13430];
assign MEM[16452] = MEM[8900] + MEM[10362];
assign MEM[16453] = MEM[8902] + MEM[11287];
assign MEM[16454] = MEM[8903] + MEM[11561];
assign MEM[16455] = MEM[8905] + MEM[13075];
assign MEM[16456] = MEM[8921] + MEM[11491];
assign MEM[16457] = MEM[8925] + MEM[9445];
assign MEM[16458] = MEM[8926] + MEM[11817];
assign MEM[16459] = MEM[8942] + MEM[11327];
assign MEM[16460] = MEM[8945] + MEM[12858];
assign MEM[16461] = MEM[8946] + MEM[10412];
assign MEM[16462] = MEM[8956] + MEM[11414];
assign MEM[16463] = MEM[8959] + MEM[9337];
assign MEM[16464] = MEM[8962] + MEM[11337];
assign MEM[16465] = MEM[8967] + MEM[14258];
assign MEM[16466] = MEM[8971] + MEM[11967];
assign MEM[16467] = MEM[8984] + MEM[12779];
assign MEM[16468] = MEM[8985] + MEM[10267];
assign MEM[16469] = MEM[8985] + MEM[10807];
assign MEM[16470] = MEM[8989] + MEM[10480];
assign MEM[16471] = MEM[8997] + MEM[10399];
assign MEM[16472] = MEM[9004] + MEM[13268];
assign MEM[16473] = MEM[9005] + MEM[11028];
assign MEM[16474] = MEM[9015] + MEM[11698];
assign MEM[16475] = MEM[9025] + MEM[9929];
assign MEM[16476] = MEM[9026] + MEM[8244];
assign MEM[16477] = MEM[9027] + MEM[13585];
assign MEM[16478] = MEM[9028] + MEM[10156];
assign MEM[16479] = MEM[9035] + MEM[11983];
assign MEM[16480] = MEM[9039] + MEM[10757];
assign MEM[16481] = MEM[9044] + MEM[9464];
assign MEM[16482] = MEM[9048] + MEM[11237];
assign MEM[16483] = MEM[9051] + MEM[10881];
assign MEM[16484] = MEM[9056] + MEM[12702];
assign MEM[16485] = MEM[9057] + MEM[11620];
assign MEM[16486] = MEM[9066] + MEM[13607];
assign MEM[16487] = MEM[9083] + MEM[11204];
assign MEM[16488] = MEM[9084] + MEM[11845];
assign MEM[16489] = MEM[9086] + MEM[13481];
assign MEM[16490] = MEM[9119] + MEM[11367];
assign MEM[16491] = MEM[9121] + MEM[11828];
assign MEM[16492] = MEM[9128] + MEM[12605];
assign MEM[16493] = MEM[9133] + MEM[10087];
assign MEM[16494] = MEM[9137] + MEM[9589];
assign MEM[16495] = MEM[9148] + MEM[10043];
assign MEM[16496] = MEM[9176] + MEM[13771];
assign MEM[16497] = MEM[9180] + MEM[11358];
assign MEM[16498] = MEM[9196] + MEM[13079];
assign MEM[16499] = MEM[9205] + MEM[11540];
assign MEM[16500] = MEM[9209] + MEM[11401];
assign MEM[16501] = MEM[9213] + MEM[11361];
assign MEM[16502] = MEM[9217] + MEM[5239];
assign MEM[16503] = MEM[9218] + MEM[10118];
assign MEM[16504] = MEM[9218] + MEM[13456];
assign MEM[16505] = MEM[9232] + MEM[9538];
assign MEM[16506] = MEM[9233] + MEM[6973];
assign MEM[16507] = MEM[9234] + MEM[12007];
assign MEM[16508] = MEM[9235] + MEM[9798];
assign MEM[16509] = MEM[9245] + MEM[11660];
assign MEM[16510] = MEM[9258] + MEM[10253];
assign MEM[16511] = MEM[9259] + MEM[10845];
assign MEM[16512] = MEM[9268] + MEM[10885];
assign MEM[16513] = MEM[9279] + MEM[9763];
assign MEM[16514] = MEM[9279] + MEM[11989];
assign MEM[16515] = MEM[9289] + MEM[11410];
assign MEM[16516] = MEM[9295] + MEM[10805];
assign MEM[16517] = MEM[9304] + MEM[10387];
assign MEM[16518] = MEM[9331] + MEM[10014];
assign MEM[16519] = MEM[9338] + MEM[11217];
assign MEM[16520] = MEM[9341] + MEM[14784];
assign MEM[16521] = MEM[9354] + MEM[10019];
assign MEM[16522] = MEM[9355] + MEM[11232];
assign MEM[16523] = MEM[9356] + MEM[14079];
assign MEM[16524] = MEM[9357] + MEM[10436];
assign MEM[16525] = MEM[9369] + MEM[9991];
assign MEM[16526] = MEM[9371] + MEM[13051];
assign MEM[16527] = MEM[9373] + MEM[12167];
assign MEM[16528] = MEM[9394] + MEM[13347];
assign MEM[16529] = MEM[9406] + MEM[11512];
assign MEM[16530] = MEM[9409] + MEM[957];
assign MEM[16531] = MEM[9413] + MEM[12423];
assign MEM[16532] = MEM[9416] + MEM[10152];
assign MEM[16533] = MEM[9419] + MEM[9695];
assign MEM[16534] = MEM[9426] + MEM[11852];
assign MEM[16535] = MEM[9428] + MEM[12241];
assign MEM[16536] = MEM[9429] + MEM[9606];
assign MEM[16537] = MEM[9448] + MEM[11640];
assign MEM[16538] = MEM[9461] + MEM[10614];
assign MEM[16539] = MEM[9471] + MEM[11226];
assign MEM[16540] = MEM[9472] + MEM[10446];
assign MEM[16541] = MEM[9480] + MEM[10355];
assign MEM[16542] = MEM[9481] + MEM[11628];
assign MEM[16543] = MEM[9483] + MEM[10003];
assign MEM[16544] = MEM[9488] + MEM[10350];
assign MEM[16545] = MEM[9492] + MEM[11451];
assign MEM[16546] = MEM[9503] + MEM[12551];
assign MEM[16547] = MEM[9508] + MEM[1671];
assign MEM[16548] = MEM[9511] + MEM[10394];
assign MEM[16549] = MEM[9516] + MEM[11400];
assign MEM[16550] = MEM[9522] + MEM[9633];
assign MEM[16551] = MEM[9527] + MEM[10499];
assign MEM[16552] = MEM[9528] + MEM[10521];
assign MEM[16553] = MEM[9533] + MEM[11376];
assign MEM[16554] = MEM[9554] + MEM[9914];
assign MEM[16555] = MEM[9557] + MEM[9867];
assign MEM[16556] = MEM[9561] + MEM[3885];
assign MEM[16557] = MEM[9565] + MEM[10607];
assign MEM[16558] = MEM[9574] + MEM[9837];
assign MEM[16559] = MEM[9576] + MEM[10967];
assign MEM[16560] = MEM[9580] + MEM[8419];
assign MEM[16561] = MEM[9583] + MEM[9906];
assign MEM[16562] = MEM[9586] + MEM[8004];
assign MEM[16563] = MEM[9587] + MEM[7042];
assign MEM[16564] = MEM[9597] + MEM[8025];
assign MEM[16565] = MEM[9602] + MEM[12415];
assign MEM[16566] = MEM[9607] + MEM[10066];
assign MEM[16567] = MEM[9609] + MEM[11503];
assign MEM[16568] = MEM[9618] + MEM[9808];
assign MEM[16569] = MEM[9624] + MEM[10806];
assign MEM[16570] = MEM[9630] + MEM[10592];
assign MEM[16571] = MEM[9637] + MEM[11214];
assign MEM[16572] = MEM[9638] + MEM[4282];
assign MEM[16573] = MEM[9645] + MEM[13688];
assign MEM[16574] = MEM[9656] + MEM[9978];
assign MEM[16575] = MEM[9664] + MEM[9742];
assign MEM[16576] = MEM[9670] + MEM[10759];
assign MEM[16577] = MEM[9673] + MEM[12934];
assign MEM[16578] = MEM[9683] + MEM[2555];
assign MEM[16579] = MEM[9692] + MEM[10694];
assign MEM[16580] = MEM[9694] + MEM[12579];
assign MEM[16581] = MEM[9700] + MEM[9903];
assign MEM[16582] = MEM[9702] + MEM[9766];
assign MEM[16583] = MEM[9712] + MEM[10371];
assign MEM[16584] = MEM[9713] + MEM[10084];
assign MEM[16585] = MEM[9727] + MEM[10352];
assign MEM[16586] = MEM[9727] + MEM[13464];
assign MEM[16587] = MEM[9730] + MEM[10646];
assign MEM[16588] = MEM[9741] + MEM[9790];
assign MEM[16589] = MEM[9744] + MEM[11514];
assign MEM[16590] = MEM[9746] + MEM[9975];
assign MEM[16591] = MEM[9748] + MEM[6706];
assign MEM[16592] = MEM[9748] + MEM[13361];
assign MEM[16593] = MEM[9758] + MEM[12642];
assign MEM[16594] = MEM[9762] + MEM[10294];
assign MEM[16595] = MEM[9763] + MEM[10581];
assign MEM[16596] = MEM[9775] + MEM[10602];
assign MEM[16597] = MEM[9782] + MEM[11618];
assign MEM[16598] = MEM[9791] + MEM[10612];
assign MEM[16599] = MEM[9803] + MEM[12896];
assign MEM[16600] = MEM[9812] + MEM[11969];
assign MEM[16601] = MEM[9813] + MEM[10323];
assign MEM[16602] = MEM[9822] + MEM[10439];
assign MEM[16603] = MEM[9822] + MEM[11377];
assign MEM[16604] = MEM[9826] + MEM[12289];
assign MEM[16605] = MEM[9838] + MEM[3029];
assign MEM[16606] = MEM[9846] + MEM[7463];
assign MEM[16607] = MEM[9847] + MEM[2309];
assign MEM[16608] = MEM[9851] + MEM[10896];
assign MEM[16609] = MEM[9869] + MEM[3845];
assign MEM[16610] = MEM[9870] + MEM[10274];
assign MEM[16611] = MEM[9873] + MEM[10160];
assign MEM[16612] = MEM[9877] + MEM[10296];
assign MEM[16613] = MEM[9877] + MEM[11611];
assign MEM[16614] = MEM[9884] + MEM[11508];
assign MEM[16615] = MEM[9891] + MEM[15211];
assign MEM[16616] = MEM[9894] + MEM[10268];
assign MEM[16617] = MEM[9896] + MEM[11707];
assign MEM[16618] = MEM[9899] + MEM[10395];
assign MEM[16619] = MEM[9904] + MEM[10196];
assign MEM[16620] = MEM[9912] + MEM[10519];
assign MEM[16621] = MEM[9920] + MEM[7455];
assign MEM[16622] = MEM[9930] + MEM[11500];
assign MEM[16623] = MEM[9932] + MEM[2059];
assign MEM[16624] = MEM[9935] + MEM[3683];
assign MEM[16625] = MEM[9937] + MEM[10107];
assign MEM[16626] = MEM[9939] + MEM[10075];
assign MEM[16627] = MEM[9943] + MEM[12009];
assign MEM[16628] = MEM[9946] + MEM[13521];
assign MEM[16629] = MEM[9949] + MEM[9123];
assign MEM[16630] = MEM[9954] + MEM[11549];
assign MEM[16631] = MEM[9967] + MEM[10925];
assign MEM[16632] = MEM[9970] + MEM[4130];
assign MEM[16633] = MEM[9981] + MEM[10146];
assign MEM[16634] = MEM[9983] + MEM[11333];
assign MEM[16635] = MEM[9987] + MEM[11588];
assign MEM[16636] = MEM[9996] + MEM[10074];
assign MEM[16637] = MEM[9997] + MEM[11282];
assign MEM[16638] = MEM[9999] + MEM[10243];
assign MEM[16639] = MEM[10004] + MEM[10481];
assign MEM[16640] = MEM[10008] + MEM[3619];
assign MEM[16641] = MEM[10009] + MEM[11350];
assign MEM[16642] = MEM[10017] + MEM[10624];
assign MEM[16643] = MEM[10030] + MEM[10429];
assign MEM[16644] = MEM[10032] + MEM[10239];
assign MEM[16645] = MEM[10033] + MEM[8396];
assign MEM[16646] = MEM[10035] + MEM[10058];
assign MEM[16647] = MEM[10037] + MEM[12614];
assign MEM[16648] = MEM[10047] + MEM[13736];
assign MEM[16649] = MEM[10063] + MEM[11735];
assign MEM[16650] = MEM[10063] + MEM[11957];
assign MEM[16651] = MEM[10068] + MEM[13349];
assign MEM[16652] = MEM[10070] + MEM[7886];
assign MEM[16653] = MEM[10093] + MEM[10365];
assign MEM[16654] = MEM[10104] + MEM[11907];
assign MEM[16655] = MEM[10105] + MEM[11222];
assign MEM[16656] = MEM[10106] + MEM[10672];
assign MEM[16657] = MEM[10109] + MEM[11454];
assign MEM[16658] = MEM[10115] + MEM[10493];
assign MEM[16659] = MEM[10119] + MEM[10202];
assign MEM[16660] = MEM[10120] + MEM[10876];
assign MEM[16661] = MEM[10120] + MEM[15477];
assign MEM[16662] = MEM[10122] + MEM[10149];
assign MEM[16663] = MEM[10127] + MEM[10494];
assign MEM[16664] = MEM[10130] + MEM[11690];
assign MEM[16665] = MEM[10133] + MEM[10697];
assign MEM[16666] = MEM[10135] + MEM[11718];
assign MEM[16667] = MEM[10150] + MEM[10263];
assign MEM[16668] = MEM[10158] + MEM[10427];
assign MEM[16669] = MEM[10159] + MEM[11964];
assign MEM[16670] = MEM[10159] + MEM[12974];
assign MEM[16671] = MEM[10161] + MEM[7648];
assign MEM[16672] = MEM[10165] + MEM[10514];
assign MEM[16673] = MEM[10167] + MEM[7964];
assign MEM[16674] = MEM[10174] + MEM[11832];
assign MEM[16675] = MEM[10183] + MEM[12783];
assign MEM[16676] = MEM[10185] + MEM[11751];
assign MEM[16677] = MEM[10185] + MEM[15360];
assign MEM[16678] = MEM[10193] + MEM[10509];
assign MEM[16679] = MEM[10195] + MEM[10289];
assign MEM[16680] = MEM[10198] + MEM[11339];
assign MEM[16681] = MEM[10199] + MEM[5861];
assign MEM[16682] = MEM[10200] + MEM[10363];
assign MEM[16683] = MEM[10205] + MEM[10723];
assign MEM[16684] = MEM[10207] + MEM[10423];
assign MEM[16685] = MEM[10219] + MEM[12221];
assign MEM[16686] = MEM[10222] + MEM[10939];
assign MEM[16687] = MEM[10224] + MEM[10977];
assign MEM[16688] = MEM[10229] + MEM[11009];
assign MEM[16689] = MEM[10231] + MEM[12054];
assign MEM[16690] = MEM[10233] + MEM[10622];
assign MEM[16691] = MEM[10234] + MEM[11138];
assign MEM[16692] = MEM[10235] + MEM[11955];
assign MEM[16693] = MEM[10240] + MEM[11420];
assign MEM[16694] = MEM[10241] + MEM[13684];
assign MEM[16695] = MEM[10242] + MEM[8588];
assign MEM[16696] = MEM[10247] + MEM[11970];
assign MEM[16697] = MEM[10254] + MEM[5518];
assign MEM[16698] = MEM[10256] + MEM[9649];
assign MEM[16699] = MEM[10261] + MEM[10542];
assign MEM[16700] = MEM[10264] + MEM[11193];
assign MEM[16701] = MEM[10266] + MEM[11719];
assign MEM[16702] = MEM[10272] + MEM[11481];
assign MEM[16703] = MEM[10273] + MEM[10838];
assign MEM[16704] = MEM[10280] + MEM[7947];
assign MEM[16705] = MEM[10280] + MEM[13173];
assign MEM[16706] = MEM[10283] + MEM[12464];
assign MEM[16707] = MEM[10283] + MEM[13138];
assign MEM[16708] = MEM[10285] + MEM[11738];
assign MEM[16709] = MEM[10286] + MEM[11729];
assign MEM[16710] = MEM[10290] + MEM[10324];
assign MEM[16711] = MEM[10299] + MEM[10326];
assign MEM[16712] = MEM[10300] + MEM[10673];
assign MEM[16713] = MEM[10303] + MEM[12639];
assign MEM[16714] = MEM[10310] + MEM[11912];
assign MEM[16715] = MEM[10316] + MEM[2397];
assign MEM[16716] = MEM[10317] + MEM[10731];
assign MEM[16717] = MEM[10320] + MEM[4237];
assign MEM[16718] = MEM[10321] + MEM[11364];
assign MEM[16719] = MEM[10322] + MEM[10670];
assign MEM[16720] = MEM[10330] + MEM[7884];
assign MEM[16721] = MEM[10332] + MEM[13812];
assign MEM[16722] = MEM[10333] + MEM[11651];
assign MEM[16723] = MEM[10334] + MEM[11304];
assign MEM[16724] = MEM[10336] + MEM[9050];
assign MEM[16725] = MEM[10337] + MEM[11303];
assign MEM[16726] = MEM[10339] + MEM[4686];
assign MEM[16727] = MEM[10341] + MEM[8610];
assign MEM[16728] = MEM[10343] + MEM[8464];
assign MEM[16729] = MEM[10346] + MEM[10588];
assign MEM[16730] = MEM[10349] + MEM[10360];
assign MEM[16731] = MEM[10353] + MEM[12040];
assign MEM[16732] = MEM[10361] + MEM[12148];
assign MEM[16733] = MEM[10366] + MEM[1331];
assign MEM[16734] = MEM[10368] + MEM[11321];
assign MEM[16735] = MEM[10370] + MEM[14594];
assign MEM[16736] = MEM[10378] + MEM[10537];
assign MEM[16737] = MEM[10381] + MEM[10398];
assign MEM[16738] = MEM[10388] + MEM[10421];
assign MEM[16739] = MEM[10389] + MEM[5799];
assign MEM[16740] = MEM[10397] + MEM[10653];
assign MEM[16741] = MEM[10400] + MEM[11959];
assign MEM[16742] = MEM[10403] + MEM[11784];
assign MEM[16743] = MEM[10405] + MEM[11435];
assign MEM[16744] = MEM[10409] + MEM[10975];
assign MEM[16745] = MEM[10410] + MEM[11310];
assign MEM[16746] = MEM[10411] + MEM[12532];
assign MEM[16747] = MEM[10413] + MEM[10871];
assign MEM[16748] = MEM[10414] + MEM[11599];
assign MEM[16749] = MEM[10416] + MEM[10649];
assign MEM[16750] = MEM[10417] + MEM[12041];
assign MEM[16751] = MEM[10418] + MEM[11178];
assign MEM[16752] = MEM[10420] + MEM[7097];
assign MEM[16753] = MEM[10422] + MEM[11419];
assign MEM[16754] = MEM[10424] + MEM[12136];
assign MEM[16755] = MEM[10425] + MEM[10658];
assign MEM[16756] = MEM[10428] + MEM[11356];
assign MEM[16757] = MEM[10431] + MEM[10488];
assign MEM[16758] = MEM[10433] + MEM[10706];
assign MEM[16759] = MEM[10434] + MEM[10872];
assign MEM[16760] = MEM[10438] + MEM[10691];
assign MEM[16761] = MEM[10441] + MEM[10837];
assign MEM[16762] = MEM[10442] + MEM[12486];
assign MEM[16763] = MEM[10443] + MEM[12012];
assign MEM[16764] = MEM[10445] + MEM[11867];
assign MEM[16765] = MEM[10447] + MEM[12132];
assign MEM[16766] = MEM[10448] + MEM[2302];
assign MEM[16767] = MEM[10450] + MEM[9859];
assign MEM[16768] = MEM[10451] + MEM[11346];
assign MEM[16769] = MEM[10453] + MEM[3179];
assign MEM[16770] = MEM[10454] + MEM[10884];
assign MEM[16771] = MEM[10455] + MEM[10955];
assign MEM[16772] = MEM[10457] + MEM[10524];
assign MEM[16773] = MEM[10459] + MEM[11498];
assign MEM[16774] = MEM[10466] + MEM[10618];
assign MEM[16775] = MEM[10471] + MEM[10921];
assign MEM[16776] = MEM[10472] + MEM[11396];
assign MEM[16777] = MEM[10473] + MEM[11626];
assign MEM[16778] = MEM[10484] + MEM[11578];
assign MEM[16779] = MEM[10486] + MEM[11776];
assign MEM[16780] = MEM[10492] + MEM[10627];
assign MEM[16781] = MEM[10495] + MEM[10822];
assign MEM[16782] = MEM[10500] + MEM[4738];
assign MEM[16783] = MEM[10500] + MEM[12151];
assign MEM[16784] = MEM[10502] + MEM[1988];
assign MEM[16785] = MEM[10510] + MEM[11649];
assign MEM[16786] = MEM[10511] + MEM[11442];
assign MEM[16787] = MEM[10512] + MEM[12033];
assign MEM[16788] = MEM[10517] + MEM[11931];
assign MEM[16789] = MEM[10518] + MEM[12883];
assign MEM[16790] = MEM[10520] + MEM[11277];
assign MEM[16791] = MEM[10522] + MEM[9339];
assign MEM[16792] = MEM[10528] + MEM[2158];
assign MEM[16793] = MEM[10532] + MEM[8086];
assign MEM[16794] = MEM[10533] + MEM[10579];
assign MEM[16795] = MEM[10538] + MEM[7441];
assign MEM[16796] = MEM[10540] + MEM[10808];
assign MEM[16797] = MEM[10541] + MEM[4382];
assign MEM[16798] = MEM[10544] + MEM[1318];
assign MEM[16799] = MEM[10546] + MEM[4446];
assign MEM[16800] = MEM[10548] + MEM[11551];
assign MEM[16801] = MEM[10550] + MEM[11563];
assign MEM[16802] = MEM[10551] + MEM[11827];
assign MEM[16803] = MEM[10552] + MEM[11627];
assign MEM[16804] = MEM[10553] + MEM[12825];
assign MEM[16805] = MEM[10557] + MEM[10563];
assign MEM[16806] = MEM[10559] + MEM[10713];
assign MEM[16807] = MEM[10568] + MEM[11436];
assign MEM[16808] = MEM[10571] + MEM[10599];
assign MEM[16809] = MEM[10572] + MEM[12018];
assign MEM[16810] = MEM[10576] + MEM[11146];
assign MEM[16811] = MEM[10577] + MEM[11253];
assign MEM[16812] = MEM[10586] + MEM[13064];
assign MEM[16813] = MEM[10590] + MEM[13292];
assign MEM[16814] = MEM[10591] + MEM[12052];
assign MEM[16815] = MEM[10595] + MEM[11866];
assign MEM[16816] = MEM[10598] + MEM[12502];
assign MEM[16817] = MEM[10600] + MEM[11554];
assign MEM[16818] = MEM[10606] + MEM[11717];
assign MEM[16819] = MEM[10608] + MEM[12032];
assign MEM[16820] = MEM[10621] + MEM[11422];
assign MEM[16821] = MEM[10628] + MEM[11051];
assign MEM[16822] = MEM[10630] + MEM[10794];
assign MEM[16823] = MEM[10639] + MEM[10887];
assign MEM[16824] = MEM[10641] + MEM[6959];
assign MEM[16825] = MEM[10644] + MEM[6445];
assign MEM[16826] = MEM[10645] + MEM[11883];
assign MEM[16827] = MEM[10647] + MEM[10633];
assign MEM[16828] = MEM[10651] + MEM[11678];
assign MEM[16829] = MEM[10655] + MEM[11111];
assign MEM[16830] = MEM[10659] + MEM[11899];
assign MEM[16831] = MEM[10663] + MEM[11538];
assign MEM[16832] = MEM[10665] + MEM[7923];
assign MEM[16833] = MEM[10669] + MEM[12251];
assign MEM[16834] = MEM[10671] + MEM[7721];
assign MEM[16835] = MEM[10676] + MEM[11968];
assign MEM[16836] = MEM[10677] + MEM[11882];
assign MEM[16837] = MEM[10678] + MEM[12123];
assign MEM[16838] = MEM[10679] + MEM[11393];
assign MEM[16839] = MEM[10680] + MEM[11323];
assign MEM[16840] = MEM[10681] + MEM[12021];
assign MEM[16841] = MEM[10684] + MEM[10764];
assign MEM[16842] = MEM[10692] + MEM[12164];
assign MEM[16843] = MEM[10695] + MEM[2332];
assign MEM[16844] = MEM[10696] + MEM[11254];
assign MEM[16845] = MEM[10700] + MEM[11365];
assign MEM[16846] = MEM[10704] + MEM[2882];
assign MEM[16847] = MEM[10707] + MEM[11288];
assign MEM[16848] = MEM[10711] + MEM[11366];
assign MEM[16849] = MEM[10712] + MEM[6914];
assign MEM[16850] = MEM[10716] + MEM[11903];
assign MEM[16851] = MEM[10718] + MEM[11168];
assign MEM[16852] = MEM[10719] + MEM[11659];
assign MEM[16853] = MEM[10720] + MEM[12515];
assign MEM[16854] = MEM[10725] + MEM[4766];
assign MEM[16855] = MEM[10730] + MEM[11372];
assign MEM[16856] = MEM[10735] + MEM[13119];
assign MEM[16857] = MEM[10738] + MEM[4710];
assign MEM[16858] = MEM[10741] + MEM[7490];
assign MEM[16859] = MEM[10749] + MEM[11846];
assign MEM[16860] = MEM[10750] + MEM[11507];
assign MEM[16861] = MEM[10753] + MEM[11453];
assign MEM[16862] = MEM[10754] + MEM[11441];
assign MEM[16863] = MEM[10767] + MEM[12030];
assign MEM[16864] = MEM[10768] + MEM[11444];
assign MEM[16865] = MEM[10771] + MEM[12658];
assign MEM[16866] = MEM[10772] + MEM[10792];
assign MEM[16867] = MEM[10773] + MEM[4998];
assign MEM[16868] = MEM[10780] + MEM[11594];
assign MEM[16869] = MEM[10781] + MEM[11709];
assign MEM[16870] = MEM[10782] + MEM[10892];
assign MEM[16871] = MEM[10784] + MEM[11689];
assign MEM[16872] = MEM[10787] + MEM[11228];
assign MEM[16873] = MEM[10793] + MEM[11787];
assign MEM[16874] = MEM[10796] + MEM[11218];
assign MEM[16875] = MEM[10802] + MEM[11736];
assign MEM[16876] = MEM[10809] + MEM[10972];
assign MEM[16877] = MEM[10820] + MEM[11731];
assign MEM[16878] = MEM[10829] + MEM[10928];
assign MEM[16879] = MEM[10830] + MEM[11961];
assign MEM[16880] = MEM[10833] + MEM[12881];
assign MEM[16881] = MEM[10834] + MEM[11161];
assign MEM[16882] = MEM[10836] + MEM[10901];
assign MEM[16883] = MEM[10844] + MEM[12072];
assign MEM[16884] = MEM[10846] + MEM[11874];
assign MEM[16885] = MEM[10848] + MEM[11375];
assign MEM[16886] = MEM[10851] + MEM[12707];
assign MEM[16887] = MEM[10853] + MEM[12081];
assign MEM[16888] = MEM[10854] + MEM[12892];
assign MEM[16889] = MEM[10855] + MEM[10797];
assign MEM[16890] = MEM[10857] + MEM[11800];
assign MEM[16891] = MEM[10858] + MEM[13158];
assign MEM[16892] = MEM[10859] + MEM[11721];
assign MEM[16893] = MEM[10860] + MEM[11195];
assign MEM[16894] = MEM[10868] + MEM[12096];
assign MEM[16895] = MEM[10880] + MEM[13089];
assign MEM[16896] = MEM[10882] + MEM[13396];
assign MEM[16897] = MEM[10891] + MEM[3382];
assign MEM[16898] = MEM[10920] + MEM[11808];
assign MEM[16899] = MEM[10930] + MEM[11389];
assign MEM[16900] = MEM[10940] + MEM[11679];
assign MEM[16901] = MEM[10942] + MEM[12422];
assign MEM[16902] = MEM[10953] + MEM[12542];
assign MEM[16903] = MEM[10961] + MEM[11884];
assign MEM[16904] = MEM[10962] + MEM[11946];
assign MEM[16905] = MEM[10963] + MEM[11695];
assign MEM[16906] = MEM[10966] + MEM[7659];
assign MEM[16907] = MEM[10968] + MEM[10812];
assign MEM[16908] = MEM[10974] + MEM[12024];
assign MEM[16909] = MEM[10979] + MEM[3731];
assign MEM[16910] = MEM[11011] + MEM[12940];
assign MEM[16911] = MEM[11016] + MEM[13494];
assign MEM[16912] = MEM[11024] + MEM[11656];
assign MEM[16913] = MEM[11035] + MEM[7576];
assign MEM[16914] = MEM[11068] + MEM[13485];
assign MEM[16915] = MEM[11074] + MEM[5133];
assign MEM[16916] = MEM[11101] + MEM[11329];
assign MEM[16917] = MEM[11116] + MEM[11666];
assign MEM[16918] = MEM[11161] + MEM[11489];
assign MEM[16919] = MEM[11162] + MEM[12509];
assign MEM[16920] = MEM[11165] + MEM[11645];
assign MEM[16921] = MEM[11166] + MEM[11893];
assign MEM[16922] = MEM[11185] + MEM[6922];
assign MEM[16923] = MEM[11192] + MEM[11466];
assign MEM[16924] = MEM[11205] + MEM[11505];
assign MEM[16925] = MEM[11210] + MEM[10810];
assign MEM[16926] = MEM[11213] + MEM[11604];
assign MEM[16927] = MEM[11231] + MEM[7379];
assign MEM[16928] = MEM[11248] + MEM[10664];
assign MEM[16929] = MEM[11261] + MEM[12846];
assign MEM[16930] = MEM[11264] + MEM[11834];
assign MEM[16931] = MEM[11275] + MEM[13909];
assign MEM[16932] = MEM[11281] + MEM[11877];
assign MEM[16933] = MEM[11296] + MEM[7369];
assign MEM[16934] = MEM[11297] + MEM[15431];
assign MEM[16935] = MEM[11305] + MEM[12437];
assign MEM[16936] = MEM[11306] + MEM[12037];
assign MEM[16937] = MEM[11315] + MEM[11368];
assign MEM[16938] = MEM[11333] + MEM[13540];
assign MEM[16939] = MEM[11347] + MEM[13650];
assign MEM[16940] = MEM[11351] + MEM[11688];
assign MEM[16941] = MEM[11354] + MEM[11586];
assign MEM[16942] = MEM[11355] + MEM[13095];
assign MEM[16943] = MEM[11355] + MEM[13339];
assign MEM[16944] = MEM[11358] + MEM[11625];
assign MEM[16945] = MEM[11360] + MEM[7025];
assign MEM[16946] = MEM[11378] + MEM[12043];
assign MEM[16947] = MEM[11379] + MEM[11571];
assign MEM[16948] = MEM[11382] + MEM[4079];
assign MEM[16949] = MEM[11384] + MEM[11591];
assign MEM[16950] = MEM[11397] + MEM[11706];
assign MEM[16951] = MEM[11398] + MEM[15094];
assign MEM[16952] = MEM[11399] + MEM[12996];
assign MEM[16953] = MEM[11405] + MEM[12441];
assign MEM[16954] = MEM[11407] + MEM[12967];
assign MEM[16955] = MEM[11409] + MEM[11474];
assign MEM[16956] = MEM[11412] + MEM[13734];
assign MEM[16957] = MEM[11413] + MEM[11107];
assign MEM[16958] = MEM[11414] + MEM[14497];
assign MEM[16959] = MEM[11416] + MEM[8314];
assign MEM[16960] = MEM[11417] + MEM[11778];
assign MEM[16961] = MEM[11421] + MEM[2372];
assign MEM[16962] = MEM[11421] + MEM[13887];
assign MEM[16963] = MEM[11429] + MEM[10440];
assign MEM[16964] = MEM[11430] + MEM[6179];
assign MEM[16965] = MEM[11432] + MEM[11546];
assign MEM[16966] = MEM[11437] + MEM[11992];
assign MEM[16967] = MEM[11438] + MEM[3627];
assign MEM[16968] = MEM[11439] + MEM[11728];
assign MEM[16969] = MEM[11439] + MEM[15191];
assign MEM[16970] = MEM[11443] + MEM[11121];
assign MEM[16971] = MEM[11448] + MEM[12616];
assign MEM[16972] = MEM[11449] + MEM[11595];
assign MEM[16973] = MEM[11450] + MEM[11668];
assign MEM[16974] = MEM[11457] + MEM[8420];
assign MEM[16975] = MEM[11458] + MEM[3303];
assign MEM[16976] = MEM[11463] + MEM[12513];
assign MEM[16977] = MEM[11467] + MEM[14310];
assign MEM[16978] = MEM[11469] + MEM[5788];
assign MEM[16979] = MEM[11471] + MEM[12175];
assign MEM[16980] = MEM[11472] + MEM[12003];
assign MEM[16981] = MEM[11475] + MEM[11539];
assign MEM[16982] = MEM[11479] + MEM[4947];
assign MEM[16983] = MEM[11480] + MEM[11781];
assign MEM[16984] = MEM[11483] + MEM[6564];
assign MEM[16985] = MEM[11485] + MEM[12234];
assign MEM[16986] = MEM[11487] + MEM[13611];
assign MEM[16987] = MEM[11489] + MEM[11685];
assign MEM[16988] = MEM[11493] + MEM[11603];
assign MEM[16989] = MEM[11495] + MEM[12000];
assign MEM[16990] = MEM[11496] + MEM[11515];
assign MEM[16991] = MEM[11504] + MEM[12107];
assign MEM[16992] = MEM[11508] + MEM[13118];
assign MEM[16993] = MEM[11510] + MEM[13180];
assign MEM[16994] = MEM[11513] + MEM[8228];
assign MEM[16995] = MEM[11514] + MEM[11788];
assign MEM[16996] = MEM[11518] + MEM[12194];
assign MEM[16997] = MEM[11525] + MEM[11682];
assign MEM[16998] = MEM[11528] + MEM[12529];
assign MEM[16999] = MEM[11530] + MEM[14023];
assign MEM[17000] = MEM[11531] + MEM[11792];
assign MEM[17001] = MEM[11532] + MEM[11564];
assign MEM[17002] = MEM[11536] + MEM[3435];
assign MEM[17003] = MEM[11537] + MEM[13187];
assign MEM[17004] = MEM[11541] + MEM[12134];
assign MEM[17005] = MEM[11542] + MEM[11632];
assign MEM[17006] = MEM[11544] + MEM[12124];
assign MEM[17007] = MEM[11553] + MEM[11658];
assign MEM[17008] = MEM[11556] + MEM[12457];
assign MEM[17009] = MEM[11562] + MEM[12095];
assign MEM[17010] = MEM[11572] + MEM[11715];
assign MEM[17011] = MEM[11575] + MEM[12093];
assign MEM[17012] = MEM[11576] + MEM[2887];
assign MEM[17013] = MEM[11580] + MEM[2482];
assign MEM[17014] = MEM[11581] + MEM[12008];
assign MEM[17015] = MEM[11584] + MEM[11704];
assign MEM[17016] = MEM[11585] + MEM[11654];
assign MEM[17017] = MEM[11587] + MEM[6055];
assign MEM[17018] = MEM[11592] + MEM[6420];
assign MEM[17019] = MEM[11596] + MEM[13787];
assign MEM[17020] = MEM[11601] + MEM[10798];
assign MEM[17021] = MEM[11602] + MEM[7844];
assign MEM[17022] = MEM[11606] + MEM[10831];
assign MEM[17023] = MEM[11607] + MEM[13579];
assign MEM[17024] = MEM[11613] + MEM[5044];
assign MEM[17025] = MEM[11614] + MEM[11951];
assign MEM[17026] = MEM[11616] + MEM[12651];
assign MEM[17027] = MEM[11617] + MEM[11793];
assign MEM[17028] = MEM[11619] + MEM[12792];
assign MEM[17029] = MEM[11621] + MEM[12025];
assign MEM[17030] = MEM[11622] + MEM[12011];
assign MEM[17031] = MEM[11623] + MEM[12625];
assign MEM[17032] = MEM[11624] + MEM[5787];
assign MEM[17033] = MEM[11629] + MEM[12545];
assign MEM[17034] = MEM[11635] + MEM[11548];
assign MEM[17035] = MEM[11636] + MEM[11819];
assign MEM[17036] = MEM[11637] + MEM[11102];
assign MEM[17037] = MEM[11639] + MEM[10819];
assign MEM[17038] = MEM[11641] + MEM[13530];
assign MEM[17039] = MEM[11643] + MEM[10958];
assign MEM[17040] = MEM[11648] + MEM[6365];
assign MEM[17041] = MEM[11653] + MEM[11045];
assign MEM[17042] = MEM[11657] + MEM[8234];
assign MEM[17043] = MEM[11661] + MEM[8424];
assign MEM[17044] = MEM[11663] + MEM[7452];
assign MEM[17045] = MEM[11664] + MEM[1931];
assign MEM[17046] = MEM[11669] + MEM[11939];
assign MEM[17047] = MEM[11671] + MEM[11744];
assign MEM[17048] = MEM[11673] + MEM[12201];
assign MEM[17049] = MEM[11674] + MEM[350];
assign MEM[17050] = MEM[11675] + MEM[7550];
assign MEM[17051] = MEM[11680] + MEM[5579];
assign MEM[17052] = MEM[11681] + MEM[8710];
assign MEM[17053] = MEM[11683] + MEM[12045];
assign MEM[17054] = MEM[11691] + MEM[11944];
assign MEM[17055] = MEM[11699] + MEM[7698];
assign MEM[17056] = MEM[11700] + MEM[11737];
assign MEM[17057] = MEM[11701] + MEM[12608];
assign MEM[17058] = MEM[11702] + MEM[12159];
assign MEM[17059] = MEM[11705] + MEM[7759];
assign MEM[17060] = MEM[11708] + MEM[11863];
assign MEM[17061] = MEM[11710] + MEM[12834];
assign MEM[17062] = MEM[11723] + MEM[13259];
assign MEM[17063] = MEM[11725] + MEM[12466];
assign MEM[17064] = MEM[11726] + MEM[8124];
assign MEM[17065] = MEM[11730] + MEM[14585];
assign MEM[17066] = MEM[11732] + MEM[12703];
assign MEM[17067] = MEM[11734] + MEM[12023];
assign MEM[17068] = MEM[11739] + MEM[12421];
assign MEM[17069] = MEM[11743] + MEM[11991];
assign MEM[17070] = MEM[11749] + MEM[12230];
assign MEM[17071] = MEM[11752] + MEM[11916];
assign MEM[17072] = MEM[11754] + MEM[8339];
assign MEM[17073] = MEM[11760] + MEM[11742];
assign MEM[17074] = MEM[11762] + MEM[12995];
assign MEM[17075] = MEM[11765] + MEM[11981];
assign MEM[17076] = MEM[11766] + MEM[10821];
assign MEM[17077] = MEM[11767] + MEM[11301];
assign MEM[17078] = MEM[11771] + MEM[9154];
assign MEM[17079] = MEM[11772] + MEM[12589];
assign MEM[17080] = MEM[11774] + MEM[12170];
assign MEM[17081] = MEM[11775] + MEM[12549];
assign MEM[17082] = MEM[11782] + MEM[12993];
assign MEM[17083] = MEM[11783] + MEM[11865];
assign MEM[17084] = MEM[11790] + MEM[12259];
assign MEM[17085] = MEM[11794] + MEM[11857];
assign MEM[17086] = MEM[11797] + MEM[13190];
assign MEM[17087] = MEM[11802] + MEM[9550];
assign MEM[17088] = MEM[11803] + MEM[14377];
assign MEM[17089] = MEM[11804] + MEM[12913];
assign MEM[17090] = MEM[11805] + MEM[5859];
assign MEM[17091] = MEM[11807] + MEM[11911];
assign MEM[17092] = MEM[11809] + MEM[11850];
assign MEM[17093] = MEM[11810] + MEM[11785];
assign MEM[17094] = MEM[11812] + MEM[12001];
assign MEM[17095] = MEM[11813] + MEM[11036];
assign MEM[17096] = MEM[11814] + MEM[11897];
assign MEM[17097] = MEM[11815] + MEM[6975];
assign MEM[17098] = MEM[11816] + MEM[12383];
assign MEM[17099] = MEM[11818] + MEM[12490];
assign MEM[17100] = MEM[11821] + MEM[12957];
assign MEM[17101] = MEM[11824] + MEM[12528];
assign MEM[17102] = MEM[11825] + MEM[10748];
assign MEM[17103] = MEM[11826] + MEM[11979];
assign MEM[17104] = MEM[11833] + MEM[7151];
assign MEM[17105] = MEM[11835] + MEM[11869];
assign MEM[17106] = MEM[11837] + MEM[14449];
assign MEM[17107] = MEM[11838] + MEM[9198];
assign MEM[17108] = MEM[11840] + MEM[5948];
assign MEM[17109] = MEM[11851] + MEM[12540];
assign MEM[17110] = MEM[11855] + MEM[12181];
assign MEM[17111] = MEM[11858] + MEM[13103];
assign MEM[17112] = MEM[11859] + MEM[13298];
assign MEM[17113] = MEM[11868] + MEM[13801];
assign MEM[17114] = MEM[11875] + MEM[13264];
assign MEM[17115] = MEM[11878] + MEM[12068];
assign MEM[17116] = MEM[11879] + MEM[14335];
assign MEM[17117] = MEM[11880] + MEM[5854];
assign MEM[17118] = MEM[11881] + MEM[12801];
assign MEM[17119] = MEM[11885] + MEM[11135];
assign MEM[17120] = MEM[11886] + MEM[12184];
assign MEM[17121] = MEM[11890] + MEM[8074];
assign MEM[17122] = MEM[11892] + MEM[10756];
assign MEM[17123] = MEM[11895] + MEM[10001];
assign MEM[17124] = MEM[11900] + MEM[12343];
assign MEM[17125] = MEM[11904] + MEM[12036];
assign MEM[17126] = MEM[11906] + MEM[12216];
assign MEM[17127] = MEM[11909] + MEM[16239];
assign MEM[17128] = MEM[11914] + MEM[12287];
assign MEM[17129] = MEM[11917] + MEM[4186];
assign MEM[17130] = MEM[11918] + MEM[12050];
assign MEM[17131] = MEM[11921] + MEM[11175];
assign MEM[17132] = MEM[11923] + MEM[12867];
assign MEM[17133] = MEM[11926] + MEM[13786];
assign MEM[17134] = MEM[11929] + MEM[13654];
assign MEM[17135] = MEM[11932] + MEM[13091];
assign MEM[17136] = MEM[11933] + MEM[13526];
assign MEM[17137] = MEM[11934] + MEM[12726];
assign MEM[17138] = MEM[11936] + MEM[12609];
assign MEM[17139] = MEM[11942] + MEM[3570];
assign MEM[17140] = MEM[11943] + MEM[12305];
assign MEM[17141] = MEM[11945] + MEM[11948];
assign MEM[17142] = MEM[11947] + MEM[8539];
assign MEM[17143] = MEM[11952] + MEM[13126];
assign MEM[17144] = MEM[11953] + MEM[12246];
assign MEM[17145] = MEM[11956] + MEM[13973];
assign MEM[17146] = MEM[11958] + MEM[12530];
assign MEM[17147] = MEM[11962] + MEM[12228];
assign MEM[17148] = MEM[11963] + MEM[11066];
assign MEM[17149] = MEM[11965] + MEM[12588];
assign MEM[17150] = MEM[11966] + MEM[8884];
assign MEM[17151] = MEM[11971] + MEM[12292];
assign MEM[17152] = MEM[11977] + MEM[13482];
assign MEM[17153] = MEM[11990] + MEM[13341];
assign MEM[17154] = MEM[11993] + MEM[13113];
assign MEM[17155] = MEM[11994] + MEM[12459];
assign MEM[17156] = MEM[11995] + MEM[8952];
assign MEM[17157] = MEM[12002] + MEM[12097];
assign MEM[17158] = MEM[12004] + MEM[719];
assign MEM[17159] = MEM[12014] + MEM[11773];
assign MEM[17160] = MEM[12019] + MEM[7142];
assign MEM[17161] = MEM[12022] + MEM[12044];
assign MEM[17162] = MEM[12026] + MEM[9156];
assign MEM[17163] = MEM[12027] + MEM[11032];
assign MEM[17164] = MEM[12028] + MEM[12378];
assign MEM[17165] = MEM[12031] + MEM[13015];
assign MEM[17166] = MEM[12034] + MEM[13600];
assign MEM[17167] = MEM[12035] + MEM[11980];
assign MEM[17168] = MEM[12038] + MEM[7235];
assign MEM[17169] = MEM[12042] + MEM[13460];
assign MEM[17170] = MEM[12047] + MEM[1766];
assign MEM[17171] = MEM[12048] + MEM[3156];
assign MEM[17172] = MEM[12051] + MEM[12714];
assign MEM[17173] = MEM[12057] + MEM[6523];
assign MEM[17174] = MEM[12058] + MEM[11777];
assign MEM[17175] = MEM[12059] + MEM[12208];
assign MEM[17176] = MEM[12061] + MEM[13243];
assign MEM[17177] = MEM[12062] + MEM[12706];
assign MEM[17178] = MEM[12063] + MEM[13717];
assign MEM[17179] = MEM[12064] + MEM[13346];
assign MEM[17180] = MEM[12069] + MEM[4156];
assign MEM[17181] = MEM[12070] + MEM[11631];
assign MEM[17182] = MEM[12071] + MEM[13738];
assign MEM[17183] = MEM[12074] + MEM[12798];
assign MEM[17184] = MEM[12090] + MEM[10478];
assign MEM[17185] = MEM[12101] + MEM[10867];
assign MEM[17186] = MEM[12105] + MEM[10778];
assign MEM[17187] = MEM[12115] + MEM[12822];
assign MEM[17188] = MEM[12122] + MEM[12753];
assign MEM[17189] = MEM[12125] + MEM[12725];
assign MEM[17190] = MEM[12127] + MEM[12229];
assign MEM[17191] = MEM[12131] + MEM[3111];
assign MEM[17192] = MEM[12135] + MEM[8554];
assign MEM[17193] = MEM[12141] + MEM[7320];
assign MEM[17194] = MEM[12155] + MEM[15025];
assign MEM[17195] = MEM[12173] + MEM[5116];
assign MEM[17196] = MEM[12176] + MEM[470];
assign MEM[17197] = MEM[12198] + MEM[12406];
assign MEM[17198] = MEM[12203] + MEM[12912];
assign MEM[17199] = MEM[12204] + MEM[12085];
assign MEM[17200] = MEM[12214] + MEM[15183];
assign MEM[17201] = MEM[12217] + MEM[13591];
assign MEM[17202] = MEM[12226] + MEM[3055];
assign MEM[17203] = MEM[12231] + MEM[13012];
assign MEM[17204] = MEM[12233] + MEM[10951];
assign MEM[17205] = MEM[12235] + MEM[12358];
assign MEM[17206] = MEM[12239] + MEM[3695];
assign MEM[17207] = MEM[12243] + MEM[12367];
assign MEM[17208] = MEM[12257] + MEM[12850];
assign MEM[17209] = MEM[12264] + MEM[8284];
assign MEM[17210] = MEM[12274] + MEM[8082];
assign MEM[17211] = MEM[12291] + MEM[11103];
assign MEM[17212] = MEM[12293] + MEM[11058];
assign MEM[17213] = MEM[12301] + MEM[12839];
assign MEM[17214] = MEM[12304] + MEM[11197];
assign MEM[17215] = MEM[12306] + MEM[15085];
assign MEM[17216] = MEM[12307] + MEM[9459];
assign MEM[17217] = MEM[12309] + MEM[13796];
assign MEM[17218] = MEM[12310] + MEM[12508];
assign MEM[17219] = MEM[12313] + MEM[12258];
assign MEM[17220] = MEM[12314] + MEM[12320];
assign MEM[17221] = MEM[12315] + MEM[14492];
assign MEM[17222] = MEM[12323] + MEM[9296];
assign MEM[17223] = MEM[12330] + MEM[12316];
assign MEM[17224] = MEM[12346] + MEM[6714];
assign MEM[17225] = MEM[12354] + MEM[12659];
assign MEM[17226] = MEM[12361] + MEM[13145];
assign MEM[17227] = MEM[12379] + MEM[13566];
assign MEM[17228] = MEM[12390] + MEM[12500];
assign MEM[17229] = MEM[12396] + MEM[14244];
assign MEM[17230] = MEM[12409] + MEM[11871];
assign MEM[17231] = MEM[12412] + MEM[13296];
assign MEM[17232] = MEM[12417] + MEM[12443];
assign MEM[17233] = MEM[12419] + MEM[13670];
assign MEM[17234] = MEM[12429] + MEM[1964];
assign MEM[17235] = MEM[12431] + MEM[13189];
assign MEM[17236] = MEM[12438] + MEM[12990];
assign MEM[17237] = MEM[12456] + MEM[3302];
assign MEM[17238] = MEM[12461] + MEM[3095];
assign MEM[17239] = MEM[12479] + MEM[12563];
assign MEM[17240] = MEM[12492] + MEM[5567];
assign MEM[17241] = MEM[12511] + MEM[4491];
assign MEM[17242] = MEM[12517] + MEM[13088];
assign MEM[17243] = MEM[12543] + MEM[12585];
assign MEM[17244] = MEM[12546] + MEM[12102];
assign MEM[17245] = MEM[12554] + MEM[12803];
assign MEM[17246] = MEM[12556] + MEM[12606];
assign MEM[17247] = MEM[12562] + MEM[6725];
assign MEM[17248] = MEM[12570] + MEM[14681];
assign MEM[17249] = MEM[12580] + MEM[12800];
assign MEM[17250] = MEM[12595] + MEM[8898];
assign MEM[17251] = MEM[12597] + MEM[12746];
assign MEM[17252] = MEM[12600] + MEM[12951];
assign MEM[17253] = MEM[12615] + MEM[12738];
assign MEM[17254] = MEM[12619] + MEM[7581];
assign MEM[17255] = MEM[12621] + MEM[12015];
assign MEM[17256] = MEM[12640] + MEM[13444];
assign MEM[17257] = MEM[12647] + MEM[6697];
assign MEM[17258] = MEM[12648] + MEM[11244];
assign MEM[17259] = MEM[12667] + MEM[8370];
assign MEM[17260] = MEM[12669] + MEM[12212];
assign MEM[17261] = MEM[12678] + MEM[13726];
assign MEM[17262] = MEM[12691] + MEM[15386];
assign MEM[17263] = MEM[12695] + MEM[12745];
assign MEM[17264] = MEM[12696] + MEM[12318];
assign MEM[17265] = MEM[12705] + MEM[12550];
assign MEM[17266] = MEM[12708] + MEM[13778];
assign MEM[17267] = MEM[12713] + MEM[10508];
assign MEM[17268] = MEM[12719] + MEM[12169];
assign MEM[17269] = MEM[12721] + MEM[13610];
assign MEM[17270] = MEM[12723] + MEM[12959];
assign MEM[17271] = MEM[12731] + MEM[12244];
assign MEM[17272] = MEM[12736] + MEM[13242];
assign MEM[17273] = MEM[12742] + MEM[5335];
assign MEM[17274] = MEM[12744] + MEM[8752];
assign MEM[17275] = MEM[12759] + MEM[12924];
assign MEM[17276] = MEM[12761] + MEM[13018];
assign MEM[17277] = MEM[12764] + MEM[11216];
assign MEM[17278] = MEM[12778] + MEM[12534];
assign MEM[17279] = MEM[12788] + MEM[13664];
assign MEM[17280] = MEM[12797] + MEM[14902];
assign MEM[17281] = MEM[12802] + MEM[13013];
assign MEM[17282] = MEM[12814] + MEM[11905];
assign MEM[17283] = MEM[12824] + MEM[12944];
assign MEM[17284] = MEM[12836] + MEM[10813];
assign MEM[17285] = MEM[12837] + MEM[4829];
assign MEM[17286] = MEM[12843] + MEM[12523];
assign MEM[17287] = MEM[12853] + MEM[7798];
assign MEM[17288] = MEM[12854] + MEM[12922];
assign MEM[17289] = MEM[12857] + MEM[12636];
assign MEM[17290] = MEM[12870] + MEM[13225];
assign MEM[17291] = MEM[12871] + MEM[13541];
assign MEM[17292] = MEM[12874] + MEM[13269];
assign MEM[17293] = MEM[12875] + MEM[12339];
assign MEM[17294] = MEM[12876] + MEM[13276];
assign MEM[17295] = MEM[12891] + MEM[12177];
assign MEM[17296] = MEM[12919] + MEM[12864];
assign MEM[17297] = MEM[12935] + MEM[13112];
assign MEM[17298] = MEM[12948] + MEM[11960];
assign MEM[17299] = MEM[12968] + MEM[13470];
assign MEM[17300] = MEM[12970] + MEM[15171];
assign MEM[17301] = MEM[12975] + MEM[9351];
assign MEM[17302] = MEM[12989] + MEM[4826];
assign MEM[17303] = MEM[12992] + MEM[12496];
assign MEM[17304] = MEM[12999] + MEM[5207];
assign MEM[17305] = MEM[13004] + MEM[12635];
assign MEM[17306] = MEM[13010] + MEM[13134];
assign MEM[17307] = MEM[13028] + MEM[12630];
assign MEM[17308] = MEM[13031] + MEM[7504];
assign MEM[17309] = MEM[13035] + MEM[13123];
assign MEM[17310] = MEM[13038] + MEM[13107];
assign MEM[17311] = MEM[13043] + MEM[10969];
assign MEM[17312] = MEM[13045] + MEM[13723];
assign MEM[17313] = MEM[13063] + MEM[2614];
assign MEM[17314] = MEM[13071] + MEM[6484];
assign MEM[17315] = MEM[13078] + MEM[11727];
assign MEM[17316] = MEM[13082] + MEM[13467];
assign MEM[17317] = MEM[13097] + MEM[14263];
assign MEM[17318] = MEM[13100] + MEM[10593];
assign MEM[17319] = MEM[13101] + MEM[4327];
assign MEM[17320] = MEM[13105] + MEM[6743];
assign MEM[17321] = MEM[13106] + MEM[9475];
assign MEM[17322] = MEM[13121] + MEM[7617];
assign MEM[17323] = MEM[13142] + MEM[11303];
assign MEM[17324] = MEM[13162] + MEM[13340];
assign MEM[17325] = MEM[13188] + MEM[1444];
assign MEM[17326] = MEM[13191] + MEM[10732];
assign MEM[17327] = MEM[13192] + MEM[13127];
assign MEM[17328] = MEM[13200] + MEM[4388];
assign MEM[17329] = MEM[13219] + MEM[13258];
assign MEM[17330] = MEM[13220] + MEM[11287];
assign MEM[17331] = MEM[13230] + MEM[7898];
assign MEM[17332] = MEM[13236] + MEM[5437];
assign MEM[17333] = MEM[13249] + MEM[11279];
assign MEM[17334] = MEM[13282] + MEM[14041];
assign MEM[17335] = MEM[13286] + MEM[6313];
assign MEM[17336] = MEM[13299] + MEM[13073];
assign MEM[17337] = MEM[13308] + MEM[14224];
assign MEM[17338] = MEM[13318] + MEM[5172];
assign MEM[17339] = MEM[13325] + MEM[13380];
assign MEM[17340] = MEM[13327] + MEM[14464];
assign MEM[17341] = MEM[13334] + MEM[7858];
assign MEM[17342] = MEM[13337] + MEM[12673];
assign MEM[17343] = MEM[13344] + MEM[13519];
assign MEM[17344] = MEM[13350] + MEM[13232];
assign MEM[17345] = MEM[13364] + MEM[12572];
assign MEM[17346] = MEM[13366] + MEM[10650];
assign MEM[17347] = MEM[13374] + MEM[13741];
assign MEM[17348] = MEM[13382] + MEM[8859];
assign MEM[17349] = MEM[13383] + MEM[12187];
assign MEM[17350] = MEM[13393] + MEM[12740];
assign MEM[17351] = MEM[13403] + MEM[13486];
assign MEM[17352] = MEM[13407] + MEM[12665];
assign MEM[17353] = MEM[13413] + MEM[5731];
assign MEM[17354] = MEM[13432] + MEM[15166];
assign MEM[17355] = MEM[13433] + MEM[12377];
assign MEM[17356] = MEM[13448] + MEM[13568];
assign MEM[17357] = MEM[13454] + MEM[12712];
assign MEM[17358] = MEM[13459] + MEM[13916];
assign MEM[17359] = MEM[13468] + MEM[14158];
assign MEM[17360] = MEM[13472] + MEM[11928];
assign MEM[17361] = MEM[13491] + MEM[10769];
assign MEM[17362] = MEM[13517] + MEM[14049];
assign MEM[17363] = MEM[13525] + MEM[12895];
assign MEM[17364] = MEM[13529] + MEM[4926];
assign MEM[17365] = MEM[13534] + MEM[4870];
assign MEM[17366] = MEM[13535] + MEM[10926];
assign MEM[17367] = MEM[13545] + MEM[14630];
assign MEM[17368] = MEM[13548] + MEM[12980];
assign MEM[17369] = MEM[13549] + MEM[12470];
assign MEM[17370] = MEM[13562] + MEM[1471];
assign MEM[17371] = MEM[13578] + MEM[14106];
assign MEM[17372] = MEM[13580] + MEM[12603];
assign MEM[17373] = MEM[13583] + MEM[5205];
assign MEM[17374] = MEM[13586] + MEM[12632];
assign MEM[17375] = MEM[13613] + MEM[13196];
assign MEM[17376] = MEM[13615] + MEM[11094];
assign MEM[17377] = MEM[13626] + MEM[7774];
assign MEM[17378] = MEM[13629] + MEM[13622];
assign MEM[17379] = MEM[13663] + MEM[13152];
assign MEM[17380] = MEM[13666] + MEM[13163];
assign MEM[17381] = MEM[13704] + MEM[8163];
assign MEM[17382] = MEM[13705] + MEM[13157];
assign MEM[17383] = MEM[13709] + MEM[6110];
assign MEM[17384] = MEM[13716] + MEM[5213];
assign MEM[17385] = MEM[13732] + MEM[7399];
assign MEM[17386] = MEM[13750] + MEM[13569];
assign MEM[17387] = MEM[13760] + MEM[13205];
assign MEM[17388] = MEM[13784] + MEM[10567];
assign MEM[17389] = MEM[13792] + MEM[5319];
assign MEM[17390] = MEM[13804] + MEM[12698];
assign MEM[17391] = MEM[13810] + MEM[12694];
assign MEM[17392] = MEM[13817] + MEM[9098];
assign MEM[17393] = MEM[14008] + MEM[10137];
assign MEM[17394] = MEM[14046] + MEM[5941];
assign MEM[17395] = MEM[14048] + MEM[10898];
assign MEM[17396] = MEM[14078] + MEM[11311];
assign MEM[17397] = MEM[14084] + MEM[12782];
assign MEM[17398] = MEM[14117] + MEM[11196];
assign MEM[17399] = MEM[14120] + MEM[13390];
assign MEM[17400] = MEM[14235] + MEM[4196];
assign MEM[17401] = MEM[14243] + MEM[13564];
assign MEM[17402] = MEM[14253] + MEM[13130];
assign MEM[17403] = MEM[14387] + MEM[6263];
assign MEM[17404] = MEM[14628] + MEM[13037];
assign MEM[17405] = MEM[14660] + MEM[11570];
assign MEM[17406] = MEM[14709] + MEM[12332];
assign MEM[17407] = MEM[14830] + MEM[8706];
assign MEM[17408] = MEM[14900] + MEM[13273];
assign MEM[17409] = MEM[14966] + MEM[13159];
assign MEM[17410] = MEM[15098] + MEM[12207];
assign MEM[17411] = MEM[15100] + MEM[14024];
assign MEM[17412] = MEM[15151] + MEM[10770];
assign MEM[17413] = MEM[15163] + MEM[13789];
assign MEM[17414] = MEM[15184] + MEM[4875];
assign MEM[17415] = MEM[15248] + MEM[2850];
assign MEM[17416] = MEM[15272] + MEM[7477];
assign MEM[17417] = MEM[15300] + MEM[12489];
assign MEM[17418] = MEM[15358] + MEM[13412];
assign MEM[17419] = MEM[15495] + MEM[13355];
assign MEM[17420] = MEM[15527] + MEM[12253];
assign MEM[17421] = MEM[15544] + MEM[13181];
assign MEM[17422] = MEM[15548] + MEM[13465];
assign MEM[17423] = MEM[15566] + MEM[15210];
assign MEM[17424] = MEM[15590] + MEM[11634];
assign MEM[17425] = MEM[15602] + MEM[11988];
assign MEM[17426] = MEM[15636] + MEM[13730];
assign MEM[17427] = MEM[15637] + MEM[17088];
assign MEM[17428] = MEM[15638] + MEM[12894];
assign MEM[17429] = MEM[15649] + MEM[12199];
assign MEM[17430] = MEM[15663] + MEM[15154];
assign MEM[17431] = MEM[15675] + MEM[14178];
assign MEM[17432] = MEM[15676] + MEM[13319];
assign MEM[17433] = MEM[15713] + MEM[13420];
assign MEM[17434] = MEM[15731] + MEM[13963];
assign MEM[17435] = MEM[15749] + MEM[13715];
assign MEM[17436] = MEM[15798] + MEM[12964];
assign MEM[17437] = MEM[15799] + MEM[13815];
assign MEM[17438] = MEM[15848] + MEM[12382];
assign MEM[17439] = MEM[15857] + MEM[14273];
assign MEM[17440] = MEM[15908] + MEM[13443];
assign MEM[17441] = MEM[15967] + MEM[12433];
assign MEM[17442] = MEM[16001] + MEM[14009];
assign MEM[17443] = MEM[16020] + MEM[13631];
assign MEM[17444] = MEM[16034] + MEM[13326];
assign MEM[17445] = MEM[16057] + MEM[12270];
assign MEM[17446] = MEM[16145] + MEM[12848];
assign MEM[17447] = MEM[16150] + MEM[12497];
assign MEM[17448] = MEM[16151] + MEM[12370];
assign MEM[17449] = MEM[16176] + MEM[13284];
assign MEM[17450] = MEM[16187] + MEM[14596];
assign MEM[17451] = MEM[16212] + MEM[14955];
assign MEM[17452] = MEM[16225] + MEM[13311];
assign MEM[17453] = MEM[16257] + MEM[15330];
assign MEM[17454] = MEM[16275] + MEM[11820];
assign MEM[17455] = MEM[16309] + MEM[13211];
assign MEM[17456] = MEM[16316] + MEM[14517];
assign MEM[17457] = MEM[16324] + MEM[12587];
assign MEM[17458] = MEM[16364] + MEM[13516];
assign MEM[17459] = MEM[16483] + MEM[12601];
assign MEM[17460] = MEM[16500] + MEM[12197];
assign MEM[17461] = MEM[16546] + MEM[15403];
assign MEM[17462] = MEM[16551] + MEM[14389];
assign MEM[17463] = MEM[16760] + MEM[13195];
assign MEM[17464] = MEM[16807] + MEM[13939];
assign MEM[17465] = MEM[16808] + MEM[13372];
assign MEM[17466] = MEM[16863] + MEM[15002];
assign MEM[17467] = MEM[16875] + MEM[15111];
assign MEM[17468] = MEM[16876] + MEM[12436];
assign MEM[17469] = MEM[16904] + MEM[13763];
assign MEM[17470] = MEM[17003] + MEM[13675];
assign MEM[17471] = MEM[17080] + MEM[13839];
assign MEM[17472] = MEM[17096] + MEM[15427];
assign MEM[17473] = MEM[17132] + MEM[13744];
assign MEM[17474] = MEM[17166] + MEM[14355];
assign MEM[17475] = MEM[17183] + MEM[13618];
assign MEM[17476] = MEM[17187] + MEM[13405];
assign MEM[17477] = MEM[17231] + MEM[14026];
assign MEM[17478] = MEM[17294] + MEM[14384];
assign MEM[17479] = MEM[5] + MEM[10932];
assign MEM[17480] = MEM[6] + MEM[6336];
assign MEM[17481] = MEM[7] + MEM[10999];
assign MEM[17482] = MEM[13] + MEM[741];
assign MEM[17483] = MEM[15] + MEM[2722];
assign MEM[17484] = MEM[21] + MEM[519];
assign MEM[17485] = MEM[22] + MEM[7498];
assign MEM[17486] = MEM[23] + MEM[9208];
assign MEM[17487] = MEM[30] + MEM[798];
assign MEM[17488] = MEM[31] + MEM[8819];
assign MEM[17489] = MEM[38] + MEM[3686];
assign MEM[17490] = MEM[45] + MEM[1438];
assign MEM[17491] = MEM[46] + MEM[1059];
assign MEM[17492] = MEM[47] + MEM[13532];
assign MEM[17493] = MEM[53] + MEM[1550];
assign MEM[17494] = MEM[54] + MEM[8563];
assign MEM[17495] = MEM[61] + MEM[5122];
assign MEM[17496] = MEM[62] + MEM[13592];
assign MEM[17497] = MEM[63] + MEM[3195];
assign MEM[17498] = MEM[69] + MEM[5125];
assign MEM[17499] = MEM[70] + MEM[1014];
assign MEM[17500] = MEM[71] + MEM[3346];
assign MEM[17501] = MEM[78] + MEM[6386];
assign MEM[17502] = MEM[79] + MEM[5135];
assign MEM[17503] = MEM[86] + MEM[11057];
assign MEM[17504] = MEM[87] + MEM[9193];
assign MEM[17505] = MEM[93] + MEM[2357];
assign MEM[17506] = MEM[95] + MEM[5396];
assign MEM[17507] = MEM[107] + MEM[3445];
assign MEM[17508] = MEM[108] + MEM[319];
assign MEM[17509] = MEM[108] + MEM[11972];
assign MEM[17510] = MEM[109] + MEM[5326];
assign MEM[17511] = MEM[116] + MEM[13090];
assign MEM[17512] = MEM[117] + MEM[8183];
assign MEM[17513] = MEM[119] + MEM[5254];
assign MEM[17514] = MEM[125] + MEM[8388];
assign MEM[17515] = MEM[127] + MEM[2637];
assign MEM[17516] = MEM[134] + MEM[12242];
assign MEM[17517] = MEM[135] + MEM[4228];
assign MEM[17518] = MEM[141] + MEM[8009];
assign MEM[17519] = MEM[143] + MEM[292];
assign MEM[17520] = MEM[149] + MEM[619];
assign MEM[17521] = MEM[150] + MEM[6165];
assign MEM[17522] = MEM[157] + MEM[2038];
assign MEM[17523] = MEM[158] + MEM[2823];
assign MEM[17524] = MEM[165] + MEM[3733];
assign MEM[17525] = MEM[167] + MEM[4917];
assign MEM[17526] = MEM[175] + MEM[3815];
assign MEM[17527] = MEM[181] + MEM[6337];
assign MEM[17528] = MEM[182] + MEM[2221];
assign MEM[17529] = MEM[183] + MEM[4767];
assign MEM[17530] = MEM[190] + MEM[2276];
assign MEM[17531] = MEM[191] + MEM[16842];
assign MEM[17532] = MEM[197] + MEM[9737];
assign MEM[17533] = MEM[198] + MEM[5974];
assign MEM[17534] = MEM[199] + MEM[9455];
assign MEM[17535] = MEM[205] + MEM[307];
assign MEM[17536] = MEM[206] + MEM[6803];
assign MEM[17537] = MEM[207] + MEM[2228];
assign MEM[17538] = MEM[213] + MEM[3827];
assign MEM[17539] = MEM[214] + MEM[2282];
assign MEM[17540] = MEM[215] + MEM[7458];
assign MEM[17541] = MEM[222] + MEM[7303];
assign MEM[17542] = MEM[223] + MEM[5023];
assign MEM[17543] = MEM[229] + MEM[14997];
assign MEM[17544] = MEM[230] + MEM[12458];
assign MEM[17545] = MEM[231] + MEM[8465];
assign MEM[17546] = MEM[237] + MEM[6463];
assign MEM[17547] = MEM[238] + MEM[2971];
assign MEM[17548] = MEM[247] + MEM[3959];
assign MEM[17549] = MEM[253] + MEM[694];
assign MEM[17550] = MEM[254] + MEM[1947];
assign MEM[17551] = MEM[255] + MEM[2322];
assign MEM[17552] = MEM[261] + MEM[355];
assign MEM[17553] = MEM[262] + MEM[7687];
assign MEM[17554] = MEM[263] + MEM[2359];
assign MEM[17555] = MEM[269] + MEM[7055];
assign MEM[17556] = MEM[270] + MEM[4227];
assign MEM[17557] = MEM[276] + MEM[3189];
assign MEM[17558] = MEM[277] + MEM[1414];
assign MEM[17559] = MEM[278] + MEM[8872];
assign MEM[17560] = MEM[279] + MEM[2893];
assign MEM[17561] = MEM[283] + MEM[6629];
assign MEM[17562] = MEM[284] + MEM[5298];
assign MEM[17563] = MEM[285] + MEM[7295];
assign MEM[17564] = MEM[286] + MEM[10914];
assign MEM[17565] = MEM[287] + MEM[14054];
assign MEM[17566] = MEM[291] + MEM[14166];
assign MEM[17567] = MEM[293] + MEM[8066];
assign MEM[17568] = MEM[294] + MEM[2068];
assign MEM[17569] = MEM[295] + MEM[9534];
assign MEM[17570] = MEM[300] + MEM[8059];
assign MEM[17571] = MEM[301] + MEM[9438];
assign MEM[17572] = MEM[303] + MEM[3454];
assign MEM[17573] = MEM[306] + MEM[4599];
assign MEM[17574] = MEM[309] + MEM[15031];
assign MEM[17575] = MEM[311] + MEM[11223];
assign MEM[17576] = MEM[315] + MEM[2556];
assign MEM[17577] = MEM[316] + MEM[2582];
assign MEM[17578] = MEM[317] + MEM[9849];
assign MEM[17579] = MEM[318] + MEM[2099];
assign MEM[17580] = MEM[323] + MEM[2007];
assign MEM[17581] = MEM[324] + MEM[11010];
assign MEM[17582] = MEM[327] + MEM[13397];
assign MEM[17583] = MEM[330] + MEM[1994];
assign MEM[17584] = MEM[331] + MEM[590];
assign MEM[17585] = MEM[332] + MEM[1722];
assign MEM[17586] = MEM[333] + MEM[9473];
assign MEM[17587] = MEM[335] + MEM[10877];
assign MEM[17588] = MEM[338] + MEM[9555];
assign MEM[17589] = MEM[339] + MEM[981];
assign MEM[17590] = MEM[341] + MEM[739];
assign MEM[17591] = MEM[343] + MEM[14996];
assign MEM[17592] = MEM[347] + MEM[5971];
assign MEM[17593] = MEM[349] + MEM[2723];
assign MEM[17594] = MEM[351] + MEM[3972];
assign MEM[17595] = MEM[354] + MEM[7217];
assign MEM[17596] = MEM[356] + MEM[13021];
assign MEM[17597] = MEM[357] + MEM[11381];
assign MEM[17598] = MEM[358] + MEM[380];
assign MEM[17599] = MEM[359] + MEM[10099];
assign MEM[17600] = MEM[363] + MEM[4684];
assign MEM[17601] = MEM[364] + MEM[13846];
assign MEM[17602] = MEM[365] + MEM[2644];
assign MEM[17603] = MEM[366] + MEM[11612];
assign MEM[17604] = MEM[370] + MEM[7746];
assign MEM[17605] = MEM[371] + MEM[5845];
assign MEM[17606] = MEM[372] + MEM[3014];
assign MEM[17607] = MEM[374] + MEM[9347];
assign MEM[17608] = MEM[375] + MEM[9752];
assign MEM[17609] = MEM[381] + MEM[1404];
assign MEM[17610] = MEM[382] + MEM[1166];
assign MEM[17611] = MEM[383] + MEM[2047];
assign MEM[17612] = MEM[391] + MEM[5462];
assign MEM[17613] = MEM[395] + MEM[12277];
assign MEM[17614] = MEM[396] + MEM[14388];
assign MEM[17615] = MEM[399] + MEM[8376];
assign MEM[17616] = MEM[403] + MEM[12688];
assign MEM[17617] = MEM[404] + MEM[12110];
assign MEM[17618] = MEM[405] + MEM[9716];
assign MEM[17619] = MEM[407] + MEM[7756];
assign MEM[17620] = MEM[411] + MEM[7933];
assign MEM[17621] = MEM[413] + MEM[2646];
assign MEM[17622] = MEM[414] + MEM[12737];
assign MEM[17623] = MEM[415] + MEM[9465];
assign MEM[17624] = MEM[422] + MEM[9734];
assign MEM[17625] = MEM[423] + MEM[4075];
assign MEM[17626] = MEM[429] + MEM[11064];
assign MEM[17627] = MEM[431] + MEM[12166];
assign MEM[17628] = MEM[437] + MEM[3510];
assign MEM[17629] = MEM[438] + MEM[6172];
assign MEM[17630] = MEM[445] + MEM[1717];
assign MEM[17631] = MEM[453] + MEM[15786];
assign MEM[17632] = MEM[455] + MEM[6652];
assign MEM[17633] = MEM[462] + MEM[3563];
assign MEM[17634] = MEM[463] + MEM[7983];
assign MEM[17635] = MEM[469] + MEM[4059];
assign MEM[17636] = MEM[471] + MEM[3525];
assign MEM[17637] = MEM[477] + MEM[5564];
assign MEM[17638] = MEM[479] + MEM[10886];
assign MEM[17639] = MEM[483] + MEM[8712];
assign MEM[17640] = MEM[484] + MEM[15964];
assign MEM[17641] = MEM[486] + MEM[5043];
assign MEM[17642] = MEM[487] + MEM[760];
assign MEM[17643] = MEM[493] + MEM[3243];
assign MEM[17644] = MEM[494] + MEM[9265];
assign MEM[17645] = MEM[495] + MEM[15364];
assign MEM[17646] = MEM[502] + MEM[3614];
assign MEM[17647] = MEM[503] + MEM[6703];
assign MEM[17648] = MEM[506] + MEM[12755];
assign MEM[17649] = MEM[508] + MEM[4212];
assign MEM[17650] = MEM[509] + MEM[7355];
assign MEM[17651] = MEM[510] + MEM[1317];
assign MEM[17652] = MEM[511] + MEM[6670];
assign MEM[17653] = MEM[515] + MEM[602];
assign MEM[17654] = MEM[517] + MEM[2495];
assign MEM[17655] = MEM[518] + MEM[6866];
assign MEM[17656] = MEM[525] + MEM[14174];
assign MEM[17657] = MEM[526] + MEM[862];
assign MEM[17658] = MEM[531] + MEM[8379];
assign MEM[17659] = MEM[533] + MEM[762];
assign MEM[17660] = MEM[534] + MEM[5346];
assign MEM[17661] = MEM[539] + MEM[12098];
assign MEM[17662] = MEM[541] + MEM[6307];
assign MEM[17663] = MEM[543] + MEM[12133];
assign MEM[17664] = MEM[547] + MEM[2670];
assign MEM[17665] = MEM[548] + MEM[4916];
assign MEM[17666] = MEM[549] + MEM[10525];
assign MEM[17667] = MEM[550] + MEM[4876];
assign MEM[17668] = MEM[554] + MEM[3799];
assign MEM[17669] = MEM[555] + MEM[10839];
assign MEM[17670] = MEM[556] + MEM[12219];
assign MEM[17671] = MEM[557] + MEM[2098];
assign MEM[17672] = MEM[558] + MEM[3166];
assign MEM[17673] = MEM[559] + MEM[3763];
assign MEM[17674] = MEM[563] + MEM[14277];
assign MEM[17675] = MEM[564] + MEM[2141];
assign MEM[17676] = MEM[565] + MEM[8954];
assign MEM[17677] = MEM[566] + MEM[7920];
assign MEM[17678] = MEM[567] + MEM[12495];
assign MEM[17679] = MEM[570] + MEM[4052];
assign MEM[17680] = MEM[572] + MEM[12010];
assign MEM[17681] = MEM[573] + MEM[4725];
assign MEM[17682] = MEM[574] + MEM[13800];
assign MEM[17683] = MEM[579] + MEM[11360];
assign MEM[17684] = MEM[581] + MEM[10742];
assign MEM[17685] = MEM[583] + MEM[9442];
assign MEM[17686] = MEM[584] + MEM[585];
assign MEM[17687] = MEM[586] + MEM[4843];
assign MEM[17688] = MEM[587] + MEM[15501];
assign MEM[17689] = MEM[589] + MEM[8302];
assign MEM[17690] = MEM[591] + MEM[6054];
assign MEM[17691] = MEM[595] + MEM[10402];
assign MEM[17692] = MEM[596] + MEM[13208];
assign MEM[17693] = MEM[597] + MEM[12689];
assign MEM[17694] = MEM[598] + MEM[6198];
assign MEM[17695] = MEM[601] + MEM[8382];
assign MEM[17696] = MEM[603] + MEM[4379];
assign MEM[17697] = MEM[604] + MEM[1522];
assign MEM[17698] = MEM[605] + MEM[7043];
assign MEM[17699] = MEM[607] + MEM[4283];
assign MEM[17700] = MEM[610] + MEM[2076];
assign MEM[17701] = MEM[611] + MEM[8711];
assign MEM[17702] = MEM[613] + MEM[5510];
assign MEM[17703] = MEM[614] + MEM[2892];
assign MEM[17704] = MEM[615] + MEM[9945];
assign MEM[17705] = MEM[618] + MEM[4717];
assign MEM[17706] = MEM[623] + MEM[13250];
assign MEM[17707] = MEM[626] + MEM[4803];
assign MEM[17708] = MEM[627] + MEM[7973];
assign MEM[17709] = MEM[628] + MEM[3396];
assign MEM[17710] = MEM[630] + MEM[7376];
assign MEM[17711] = MEM[631] + MEM[15047];
assign MEM[17712] = MEM[634] + MEM[14161];
assign MEM[17713] = MEM[635] + MEM[5228];
assign MEM[17714] = MEM[636] + MEM[10615];
assign MEM[17715] = MEM[637] + MEM[3965];
assign MEM[17716] = MEM[644] + MEM[2316];
assign MEM[17717] = MEM[645] + MEM[9464];
assign MEM[17718] = MEM[651] + MEM[12308];
assign MEM[17719] = MEM[653] + MEM[13291];
assign MEM[17720] = MEM[654] + MEM[9294];
assign MEM[17721] = MEM[661] + MEM[3790];
assign MEM[17722] = MEM[662] + MEM[2351];
assign MEM[17723] = MEM[669] + MEM[9592];
assign MEM[17724] = MEM[670] + MEM[16168];
assign MEM[17725] = MEM[671] + MEM[1523];
assign MEM[17726] = MEM[677] + MEM[4380];
assign MEM[17727] = MEM[678] + MEM[12049];
assign MEM[17728] = MEM[679] + MEM[4895];
assign MEM[17729] = MEM[685] + MEM[4557];
assign MEM[17730] = MEM[686] + MEM[10549];
assign MEM[17731] = MEM[693] + MEM[10929];
assign MEM[17732] = MEM[695] + MEM[1109];
assign MEM[17733] = MEM[702] + MEM[934];
assign MEM[17734] = MEM[709] + MEM[1934];
assign MEM[17735] = MEM[710] + MEM[1063];
assign MEM[17736] = MEM[711] + MEM[3221];
assign MEM[17737] = MEM[715] + MEM[7340];
assign MEM[17738] = MEM[716] + MEM[1150];
assign MEM[17739] = MEM[717] + MEM[13676];
assign MEM[17740] = MEM[724] + MEM[7153];
assign MEM[17741] = MEM[725] + MEM[2362];
assign MEM[17742] = MEM[731] + MEM[10637];
assign MEM[17743] = MEM[732] + MEM[9440];
assign MEM[17744] = MEM[734] + MEM[11633];
assign MEM[17745] = MEM[738] + MEM[6729];
assign MEM[17746] = MEM[740] + MEM[8185];
assign MEM[17747] = MEM[745] + MEM[11720];
assign MEM[17748] = MEM[746] + MEM[2307];
assign MEM[17749] = MEM[747] + MEM[1021];
assign MEM[17750] = MEM[748] + MEM[10516];
assign MEM[17751] = MEM[749] + MEM[11308];
assign MEM[17752] = MEM[750] + MEM[9379];
assign MEM[17753] = MEM[751] + MEM[5075];
assign MEM[17754] = MEM[755] + MEM[5938];
assign MEM[17755] = MEM[756] + MEM[3738];
assign MEM[17756] = MEM[757] + MEM[9936];
assign MEM[17757] = MEM[758] + MEM[5276];
assign MEM[17758] = MEM[761] + MEM[5413];
assign MEM[17759] = MEM[763] + MEM[2748];
assign MEM[17760] = MEM[765] + MEM[5815];
assign MEM[17761] = MEM[767] + MEM[9785];
assign MEM[17762] = MEM[770] + MEM[11887];
assign MEM[17763] = MEM[771] + MEM[7859];
assign MEM[17764] = MEM[773] + MEM[5523];
assign MEM[17765] = MEM[775] + MEM[11998];
assign MEM[17766] = MEM[776] + MEM[11494];
assign MEM[17767] = MEM[778] + MEM[11235];
assign MEM[17768] = MEM[781] + MEM[10101];
assign MEM[17769] = MEM[782] + MEM[14345];
assign MEM[17770] = MEM[783] + MEM[1125];
assign MEM[17771] = MEM[787] + MEM[2142];
assign MEM[17772] = MEM[788] + MEM[7864];
assign MEM[17773] = MEM[789] + MEM[5363];
assign MEM[17774] = MEM[790] + MEM[8081];
assign MEM[17775] = MEM[791] + MEM[6953];
assign MEM[17776] = MEM[795] + MEM[12147];
assign MEM[17777] = MEM[796] + MEM[6433];
assign MEM[17778] = MEM[797] + MEM[2974];
assign MEM[17779] = MEM[799] + MEM[10402];
assign MEM[17780] = MEM[800] + MEM[5574];
assign MEM[17781] = MEM[802] + MEM[10209];
assign MEM[17782] = MEM[803] + MEM[12340];
assign MEM[17783] = MEM[805] + MEM[1958];
assign MEM[17784] = MEM[806] + MEM[2327];
assign MEM[17785] = MEM[807] + MEM[11047];
assign MEM[17786] = MEM[812] + MEM[2869];
assign MEM[17787] = MEM[813] + MEM[10736];
assign MEM[17788] = MEM[814] + MEM[12260];
assign MEM[17789] = MEM[815] + MEM[5534];
assign MEM[17790] = MEM[819] + MEM[5927];
assign MEM[17791] = MEM[820] + MEM[8912];
assign MEM[17792] = MEM[822] + MEM[2335];
assign MEM[17793] = MEM[823] + MEM[3317];
assign MEM[17794] = MEM[826] + MEM[17042];
assign MEM[17795] = MEM[827] + MEM[13395];
assign MEM[17796] = MEM[828] + MEM[2051];
assign MEM[17797] = MEM[829] + MEM[2714];
assign MEM[17798] = MEM[830] + MEM[12835];
assign MEM[17799] = MEM[831] + MEM[1028];
assign MEM[17800] = MEM[834] + MEM[5676];
assign MEM[17801] = MEM[837] + MEM[11080];
assign MEM[17802] = MEM[839] + MEM[14272];
assign MEM[17803] = MEM[844] + MEM[8560];
assign MEM[17804] = MEM[845] + MEM[17435];
assign MEM[17805] = MEM[846] + MEM[11291];
assign MEM[17806] = MEM[851] + MEM[3460];
assign MEM[17807] = MEM[853] + MEM[6005];
assign MEM[17808] = MEM[854] + MEM[4967];
assign MEM[17809] = MEM[855] + MEM[8540];
assign MEM[17810] = MEM[859] + MEM[3764];
assign MEM[17811] = MEM[860] + MEM[1463];
assign MEM[17812] = MEM[861] + MEM[12512];
assign MEM[17813] = MEM[863] + MEM[1743];
assign MEM[17814] = MEM[866] + MEM[8880];
assign MEM[17815] = MEM[869] + MEM[14855];
assign MEM[17816] = MEM[874] + MEM[2117];
assign MEM[17817] = MEM[875] + MEM[2710];
assign MEM[17818] = MEM[877] + MEM[11119];
assign MEM[17819] = MEM[878] + MEM[4732];
assign MEM[17820] = MEM[879] + MEM[8860];
assign MEM[17821] = MEM[885] + MEM[2565];
assign MEM[17822] = MEM[886] + MEM[3039];
assign MEM[17823] = MEM[893] + MEM[12142];
assign MEM[17824] = MEM[894] + MEM[13484];
assign MEM[17825] = MEM[901] + MEM[9582];
assign MEM[17826] = MEM[902] + MEM[9892];
assign MEM[17827] = MEM[903] + MEM[5367];
assign MEM[17828] = MEM[909] + MEM[8141];
assign MEM[17829] = MEM[911] + MEM[1644];
assign MEM[17830] = MEM[919] + MEM[3839];
assign MEM[17831] = MEM[925] + MEM[11020];
assign MEM[17832] = MEM[927] + MEM[3866];
assign MEM[17833] = MEM[930] + MEM[4515];
assign MEM[17834] = MEM[931] + MEM[2293];
assign MEM[17835] = MEM[932] + MEM[4565];
assign MEM[17836] = MEM[933] + MEM[13034];
assign MEM[17837] = MEM[935] + MEM[13968];
assign MEM[17838] = MEM[938] + MEM[12006];
assign MEM[17839] = MEM[940] + MEM[7210];
assign MEM[17840] = MEM[941] + MEM[3082];
assign MEM[17841] = MEM[946] + MEM[5452];
assign MEM[17842] = MEM[947] + MEM[1972];
assign MEM[17843] = MEM[949] + MEM[2656];
assign MEM[17844] = MEM[950] + MEM[1260];
assign MEM[17845] = MEM[951] + MEM[9319];
assign MEM[17846] = MEM[954] + MEM[9139];
assign MEM[17847] = MEM[956] + MEM[1516];
assign MEM[17848] = MEM[958] + MEM[2108];
assign MEM[17849] = MEM[962] + MEM[13348];
assign MEM[17850] = MEM[963] + MEM[6486];
assign MEM[17851] = MEM[964] + MEM[7621];
assign MEM[17852] = MEM[965] + MEM[3018];
assign MEM[17853] = MEM[966] + MEM[10913];
assign MEM[17854] = MEM[967] + MEM[12962];
assign MEM[17855] = MEM[970] + MEM[1687];
assign MEM[17856] = MEM[971] + MEM[11894];
assign MEM[17857] = MEM[972] + MEM[2388];
assign MEM[17858] = MEM[974] + MEM[5509];
assign MEM[17859] = MEM[975] + MEM[16945];
assign MEM[17860] = MEM[978] + MEM[5268];
assign MEM[17861] = MEM[979] + MEM[13785];
assign MEM[17862] = MEM[983] + MEM[8045];
assign MEM[17863] = MEM[986] + MEM[3870];
assign MEM[17864] = MEM[987] + MEM[4541];
assign MEM[17865] = MEM[988] + MEM[13512];
assign MEM[17866] = MEM[989] + MEM[8006];
assign MEM[17867] = MEM[991] + MEM[2223];
assign MEM[17868] = MEM[994] + MEM[1175];
assign MEM[17869] = MEM[1004] + MEM[8996];
assign MEM[17870] = MEM[1006] + MEM[15650];
assign MEM[17871] = MEM[1007] + MEM[5117];
assign MEM[17872] = MEM[1011] + MEM[15446];
assign MEM[17873] = MEM[1012] + MEM[4548];
assign MEM[17874] = MEM[1013] + MEM[7658];
assign MEM[17875] = MEM[1015] + MEM[2981];
assign MEM[17876] = MEM[1019] + MEM[12861];
assign MEM[17877] = MEM[1020] + MEM[1242];
assign MEM[17878] = MEM[1022] + MEM[8736];
assign MEM[17879] = MEM[1023] + MEM[4347];
assign MEM[17880] = MEM[1026] + MEM[2701];
assign MEM[17881] = MEM[1027] + MEM[2365];
assign MEM[17882] = MEM[1030] + MEM[6182];
assign MEM[17883] = MEM[1031] + MEM[3868];
assign MEM[17884] = MEM[1034] + MEM[3872];
assign MEM[17885] = MEM[1037] + MEM[11557];
assign MEM[17886] = MEM[1038] + MEM[9480];
assign MEM[17887] = MEM[1043] + MEM[5005];
assign MEM[17888] = MEM[1044] + MEM[7218];
assign MEM[17889] = MEM[1045] + MEM[1363];
assign MEM[17890] = MEM[1046] + MEM[11401];
assign MEM[17891] = MEM[1050] + MEM[12395];
assign MEM[17892] = MEM[1051] + MEM[10497];
assign MEM[17893] = MEM[1055] + MEM[11692];
assign MEM[17894] = MEM[1058] + MEM[3562];
assign MEM[17895] = MEM[1060] + MEM[7006];
assign MEM[17896] = MEM[1061] + MEM[3522];
assign MEM[17897] = MEM[1062] + MEM[4651];
assign MEM[17898] = MEM[1067] + MEM[5786];
assign MEM[17899] = MEM[1068] + MEM[3923];
assign MEM[17900] = MEM[1069] + MEM[4676];
assign MEM[17901] = MEM[1071] + MEM[16350];
assign MEM[17902] = MEM[1074] + MEM[3063];
assign MEM[17903] = MEM[1075] + MEM[2934];
assign MEM[17904] = MEM[1076] + MEM[1278];
assign MEM[17905] = MEM[1078] + MEM[8379];
assign MEM[17906] = MEM[1082] + MEM[5500];
assign MEM[17907] = MEM[1083] + MEM[10804];
assign MEM[17908] = MEM[1085] + MEM[10570];
assign MEM[17909] = MEM[1086] + MEM[5606];
assign MEM[17910] = MEM[1090] + MEM[13596];
assign MEM[17911] = MEM[1092] + MEM[8095];
assign MEM[17912] = MEM[1093] + MEM[11370];
assign MEM[17913] = MEM[1094] + MEM[1251];
assign MEM[17914] = MEM[1095] + MEM[1276];
assign MEM[17915] = MEM[1099] + MEM[4994];
assign MEM[17916] = MEM[1101] + MEM[3831];
assign MEM[17917] = MEM[1102] + MEM[3670];
assign MEM[17918] = MEM[1103] + MEM[11042];
assign MEM[17919] = MEM[1107] + MEM[2092];
assign MEM[17920] = MEM[1110] + MEM[8075];
assign MEM[17921] = MEM[1111] + MEM[7607];
assign MEM[17922] = MEM[1119] + MEM[5253];
assign MEM[17923] = MEM[1126] + MEM[12303];
assign MEM[17924] = MEM[1133] + MEM[3391];
assign MEM[17925] = MEM[1134] + MEM[3523];
assign MEM[17926] = MEM[1135] + MEM[12670];
assign MEM[17927] = MEM[1141] + MEM[6715];
assign MEM[17928] = MEM[1142] + MEM[4372];
assign MEM[17929] = MEM[1143] + MEM[5499];
assign MEM[17930] = MEM[1147] + MEM[10422];
assign MEM[17931] = MEM[1148] + MEM[2612];
assign MEM[17932] = MEM[1149] + MEM[15988];
assign MEM[17933] = MEM[1151] + MEM[10449];
assign MEM[17934] = MEM[1154] + MEM[8833];
assign MEM[17935] = MEM[1155] + MEM[4662];
assign MEM[17936] = MEM[1156] + MEM[5674];
assign MEM[17937] = MEM[1158] + MEM[4950];
assign MEM[17938] = MEM[1162] + MEM[4605];
assign MEM[17939] = MEM[1164] + MEM[4038];
assign MEM[17940] = MEM[1165] + MEM[8437];
assign MEM[17941] = MEM[1167] + MEM[16272];
assign MEM[17942] = MEM[1170] + MEM[12076];
assign MEM[17943] = MEM[1171] + MEM[11552];
assign MEM[17944] = MEM[1172] + MEM[12945];
assign MEM[17945] = MEM[1178] + MEM[5923];
assign MEM[17946] = MEM[1179] + MEM[12223];
assign MEM[17947] = MEM[1190] + MEM[2274];
assign MEM[17948] = MEM[1191] + MEM[5195];
assign MEM[17949] = MEM[1195] + MEM[9249];
assign MEM[17950] = MEM[1197] + MEM[11283];
assign MEM[17951] = MEM[1199] + MEM[10852];
assign MEM[17952] = MEM[1202] + MEM[13769];
assign MEM[17953] = MEM[1204] + MEM[13806];
assign MEM[17954] = MEM[1205] + MEM[4399];
assign MEM[17955] = MEM[1206] + MEM[9493];
assign MEM[17956] = MEM[1211] + MEM[8294];
assign MEM[17957] = MEM[1212] + MEM[2820];
assign MEM[17958] = MEM[1213] + MEM[3474];
assign MEM[17959] = MEM[1214] + MEM[2506];
assign MEM[17960] = MEM[1215] + MEM[4117];
assign MEM[17961] = MEM[1218] + MEM[6302];
assign MEM[17962] = MEM[1223] + MEM[6287];
assign MEM[17963] = MEM[1227] + MEM[8844];
assign MEM[17964] = MEM[1228] + MEM[8019];
assign MEM[17965] = MEM[1229] + MEM[15409];
assign MEM[17966] = MEM[1235] + MEM[10597];
assign MEM[17967] = MEM[1236] + MEM[3103];
assign MEM[17968] = MEM[1238] + MEM[4412];
assign MEM[17969] = MEM[1239] + MEM[4819];
assign MEM[17970] = MEM[1246] + MEM[8574];
assign MEM[17971] = MEM[1252] + MEM[9613];
assign MEM[17972] = MEM[1253] + MEM[2811];
assign MEM[17973] = MEM[1255] + MEM[1940];
assign MEM[17974] = MEM[1259] + MEM[6492];
assign MEM[17975] = MEM[1261] + MEM[10631];
assign MEM[17976] = MEM[1262] + MEM[11072];
assign MEM[17977] = MEM[1263] + MEM[4471];
assign MEM[17978] = MEM[1266] + MEM[12252];
assign MEM[17979] = MEM[1268] + MEM[12180];
assign MEM[17980] = MEM[1269] + MEM[10648];
assign MEM[17981] = MEM[1270] + MEM[5311];
assign MEM[17982] = MEM[1271] + MEM[7483];
assign MEM[17983] = MEM[1277] + MEM[1399];
assign MEM[17984] = MEM[1283] + MEM[6753];
assign MEM[17985] = MEM[1285] + MEM[12955];
assign MEM[17986] = MEM[1286] + MEM[4019];
assign MEM[17987] = MEM[1287] + MEM[4476];
assign MEM[17988] = MEM[1291] + MEM[11742];
assign MEM[17989] = MEM[1292] + MEM[5429];
assign MEM[17990] = MEM[1293] + MEM[7876];
assign MEM[17991] = MEM[1294] + MEM[2767];
assign MEM[17992] = MEM[1295] + MEM[2078];
assign MEM[17993] = MEM[1298] + MEM[1332];
assign MEM[17994] = MEM[1300] + MEM[3237];
assign MEM[17995] = MEM[1302] + MEM[4746];
assign MEM[17996] = MEM[1303] + MEM[7633];
assign MEM[17997] = MEM[1306] + MEM[7258];
assign MEM[17998] = MEM[1307] + MEM[6744];
assign MEM[17999] = MEM[1308] + MEM[4971];
assign MEM[18000] = MEM[1309] + MEM[1507];
assign MEM[18001] = MEM[1310] + MEM[2445];
assign MEM[18002] = MEM[1311] + MEM[12487];
assign MEM[18003] = MEM[1315] + MEM[15215];
assign MEM[18004] = MEM[1319] + MEM[2350];
assign MEM[18005] = MEM[1322] + MEM[5829];
assign MEM[18006] = MEM[1323] + MEM[6428];
assign MEM[18007] = MEM[1324] + MEM[6211];
assign MEM[18008] = MEM[1325] + MEM[13466];
assign MEM[18009] = MEM[1326] + MEM[2950];
assign MEM[18010] = MEM[1327] + MEM[1349];
assign MEM[18011] = MEM[1330] + MEM[6901];
assign MEM[18012] = MEM[1335] + MEM[2525];
assign MEM[18013] = MEM[1342] + MEM[2183];
assign MEM[18014] = MEM[1351] + MEM[14958];
assign MEM[18015] = MEM[1357] + MEM[5115];
assign MEM[18016] = MEM[1358] + MEM[3611];
assign MEM[18017] = MEM[1359] + MEM[2107];
assign MEM[18018] = MEM[1367] + MEM[7275];
assign MEM[18019] = MEM[1370] + MEM[10511];
assign MEM[18020] = MEM[1371] + MEM[1900];
assign MEM[18021] = MEM[1372] + MEM[11437];
assign MEM[18022] = MEM[1374] + MEM[10982];
assign MEM[18023] = MEM[1375] + MEM[6878];
assign MEM[18024] = MEM[1378] + MEM[2278];
assign MEM[18025] = MEM[1379] + MEM[6612];
assign MEM[18026] = MEM[1380] + MEM[1779];
assign MEM[18027] = MEM[1381] + MEM[8797];
assign MEM[18028] = MEM[1386] + MEM[7744];
assign MEM[18029] = MEM[1387] + MEM[8512];
assign MEM[18030] = MEM[1388] + MEM[5476];
assign MEM[18031] = MEM[1389] + MEM[4655];
assign MEM[18032] = MEM[1390] + MEM[3823];
assign MEM[18033] = MEM[1394] + MEM[9779];
assign MEM[18034] = MEM[1396] + MEM[5373];
assign MEM[18035] = MEM[1397] + MEM[2485];
assign MEM[18036] = MEM[1398] + MEM[8523];
assign MEM[18037] = MEM[1402] + MEM[5566];
assign MEM[18038] = MEM[1403] + MEM[3903];
assign MEM[18039] = MEM[1405] + MEM[4661];
assign MEM[18040] = MEM[1410] + MEM[5886];
assign MEM[18041] = MEM[1419] + MEM[9231];
assign MEM[18042] = MEM[1421] + MEM[6584];
assign MEM[18043] = MEM[1422] + MEM[3899];
assign MEM[18044] = MEM[1423] + MEM[5997];
assign MEM[18045] = MEM[1426] + MEM[9666];
assign MEM[18046] = MEM[1427] + MEM[7972];
assign MEM[18047] = MEM[1428] + MEM[5822];
assign MEM[18048] = MEM[1429] + MEM[8517];
assign MEM[18049] = MEM[1437] + MEM[5389];
assign MEM[18050] = MEM[1439] + MEM[8961];
assign MEM[18051] = MEM[1445] + MEM[3782];
assign MEM[18052] = MEM[1446] + MEM[4060];
assign MEM[18053] = MEM[1453] + MEM[4757];
assign MEM[18054] = MEM[1454] + MEM[13141];
assign MEM[18055] = MEM[1455] + MEM[8647];
assign MEM[18056] = MEM[1458] + MEM[5469];
assign MEM[18057] = MEM[1459] + MEM[4226];
assign MEM[18058] = MEM[1461] + MEM[1594];
assign MEM[18059] = MEM[1462] + MEM[6368];
assign MEM[18060] = MEM[1466] + MEM[12077];
assign MEM[18061] = MEM[1467] + MEM[3915];
assign MEM[18062] = MEM[1470] + MEM[12245];
assign MEM[18063] = MEM[1477] + MEM[3780];
assign MEM[18064] = MEM[1478] + MEM[1812];
assign MEM[18065] = MEM[1479] + MEM[9584];
assign MEM[18066] = MEM[1483] + MEM[5366];
assign MEM[18067] = MEM[1485] + MEM[13199];
assign MEM[18068] = MEM[1487] + MEM[12602];
assign MEM[18069] = MEM[1491] + MEM[11861];
assign MEM[18070] = MEM[1501] + MEM[2895];
assign MEM[18071] = MEM[1503] + MEM[2236];
assign MEM[18072] = MEM[1506] + MEM[8756];
assign MEM[18073] = MEM[1508] + MEM[16426];
assign MEM[18074] = MEM[1510] + MEM[2798];
assign MEM[18075] = MEM[1511] + MEM[4007];
assign MEM[18076] = MEM[1514] + MEM[9545];
assign MEM[18077] = MEM[1517] + MEM[5178];
assign MEM[18078] = MEM[1518] + MEM[3579];
assign MEM[18079] = MEM[1523] + MEM[3069];
assign MEM[18080] = MEM[1527] + MEM[4501];
assign MEM[18081] = MEM[1528] + MEM[6162];
assign MEM[18082] = MEM[1531] + MEM[10976];
assign MEM[18083] = MEM[1532] + MEM[5191];
assign MEM[18084] = MEM[1533] + MEM[5245];
assign MEM[18085] = MEM[1534] + MEM[6123];
assign MEM[18086] = MEM[1535] + MEM[12586];
assign MEM[18087] = MEM[1540] + MEM[7305];
assign MEM[18088] = MEM[1542] + MEM[16819];
assign MEM[18089] = MEM[1543] + MEM[8630];
assign MEM[18090] = MEM[1546] + MEM[15359];
assign MEM[18091] = MEM[1547] + MEM[15140];
assign MEM[18092] = MEM[1551] + MEM[9497];
assign MEM[18093] = MEM[1554] + MEM[13825];
assign MEM[18094] = MEM[1555] + MEM[14203];
assign MEM[18095] = MEM[1556] + MEM[13772];
assign MEM[18096] = MEM[1558] + MEM[1862];
assign MEM[18097] = MEM[1559] + MEM[5996];
assign MEM[18098] = MEM[1563] + MEM[7940];
assign MEM[18099] = MEM[1564] + MEM[8402];
assign MEM[18100] = MEM[1566] + MEM[3867];
assign MEM[18101] = MEM[1573] + MEM[2627];
assign MEM[18102] = MEM[1574] + MEM[7987];
assign MEM[18103] = MEM[1578] + MEM[6011];
assign MEM[18104] = MEM[1580] + MEM[14891];
assign MEM[18105] = MEM[1581] + MEM[10862];
assign MEM[18106] = MEM[1582] + MEM[5757];
assign MEM[18107] = MEM[1583] + MEM[6300];
assign MEM[18108] = MEM[1587] + MEM[8763];
assign MEM[18109] = MEM[1588] + MEM[10501];
assign MEM[18110] = MEM[1589] + MEM[12535];
assign MEM[18111] = MEM[1590] + MEM[5989];
assign MEM[18112] = MEM[1591] + MEM[5765];
assign MEM[18113] = MEM[1596] + MEM[13143];
assign MEM[18114] = MEM[1598] + MEM[8155];
assign MEM[18115] = MEM[1599] + MEM[11672];
assign MEM[18116] = MEM[1602] + MEM[8667];
assign MEM[18117] = MEM[1604] + MEM[5767];
assign MEM[18118] = MEM[1605] + MEM[10060];
assign MEM[18119] = MEM[1607] + MEM[2460];
assign MEM[18120] = MEM[1610] + MEM[12449];
assign MEM[18121] = MEM[1611] + MEM[16276];
assign MEM[18122] = MEM[1612] + MEM[5934];
assign MEM[18123] = MEM[1613] + MEM[16598];
assign MEM[18124] = MEM[1614] + MEM[8901];
assign MEM[18125] = MEM[1619] + MEM[12521];
assign MEM[18126] = MEM[1621] + MEM[2563];
assign MEM[18127] = MEM[1622] + MEM[8600];
assign MEM[18128] = MEM[1623] + MEM[10919];
assign MEM[18129] = MEM[1626] + MEM[2717];
assign MEM[18130] = MEM[1627] + MEM[1876];
assign MEM[18131] = MEM[1628] + MEM[2866];
assign MEM[18132] = MEM[1629] + MEM[10464];
assign MEM[18133] = MEM[1630] + MEM[6170];
assign MEM[18134] = MEM[1634] + MEM[7445];
assign MEM[18135] = MEM[1635] + MEM[8014];
assign MEM[18136] = MEM[1636] + MEM[2493];
assign MEM[18137] = MEM[1638] + MEM[3707];
assign MEM[18138] = MEM[1639] + MEM[2301];
assign MEM[18139] = MEM[1645] + MEM[5339];
assign MEM[18140] = MEM[1646] + MEM[4972];
assign MEM[18141] = MEM[1647] + MEM[10814];
assign MEM[18142] = MEM[1650] + MEM[7888];
assign MEM[18143] = MEM[1651] + MEM[12205];
assign MEM[18144] = MEM[1652] + MEM[1948];
assign MEM[18145] = MEM[1653] + MEM[6402];
assign MEM[18146] = MEM[1659] + MEM[10949];
assign MEM[18147] = MEM[1660] + MEM[6512];
assign MEM[18148] = MEM[1661] + MEM[5890];
assign MEM[18149] = MEM[1663] + MEM[15070];
assign MEM[18150] = MEM[1667] + MEM[5299];
assign MEM[18151] = MEM[1668] + MEM[4780];
assign MEM[18152] = MEM[1676] + MEM[7414];
assign MEM[18153] = MEM[1678] + MEM[10323];
assign MEM[18154] = MEM[1679] + MEM[11930];
assign MEM[18155] = MEM[1682] + MEM[10984];
assign MEM[18156] = MEM[1683] + MEM[2222];
assign MEM[18157] = MEM[1684] + MEM[12256];
assign MEM[18158] = MEM[1685] + MEM[11896];
assign MEM[18159] = MEM[1686] + MEM[7205];
assign MEM[18160] = MEM[1690] + MEM[12997];
assign MEM[18161] = MEM[1691] + MEM[2843];
assign MEM[18162] = MEM[1693] + MEM[3786];
assign MEM[18163] = MEM[1694] + MEM[9513];
assign MEM[18164] = MEM[1695] + MEM[12961];
assign MEM[18165] = MEM[1703] + MEM[6992];
assign MEM[18166] = MEM[1707] + MEM[8605];
assign MEM[18167] = MEM[1709] + MEM[4335];
assign MEM[18168] = MEM[1710] + MEM[3668];
assign MEM[18169] = MEM[1711] + MEM[2275];
assign MEM[18170] = MEM[1715] + MEM[5703];
assign MEM[18171] = MEM[1716] + MEM[2229];
assign MEM[18172] = MEM[1718] + MEM[5679];
assign MEM[18173] = MEM[1719] + MEM[12849];
assign MEM[18174] = MEM[1723] + MEM[6378];
assign MEM[18175] = MEM[1727] + MEM[12290];
assign MEM[18176] = MEM[1730] + MEM[6012];
assign MEM[18177] = MEM[1731] + MEM[11909];
assign MEM[18178] = MEM[1732] + MEM[10248];
assign MEM[18179] = MEM[1733] + MEM[4140];
assign MEM[18180] = MEM[1734] + MEM[5495];
assign MEM[18181] = MEM[1736] + MEM[14242];
assign MEM[18182] = MEM[1739] + MEM[7453];
assign MEM[18183] = MEM[1740] + MEM[1742];
assign MEM[18184] = MEM[1746] + MEM[4341];
assign MEM[18185] = MEM[1747] + MEM[10747];
assign MEM[18186] = MEM[1748] + MEM[6117];
assign MEM[18187] = MEM[1751] + MEM[2799];
assign MEM[18188] = MEM[1756] + MEM[5069];
assign MEM[18189] = MEM[1757] + MEM[9383];
assign MEM[18190] = MEM[1758] + MEM[12209];
assign MEM[18191] = MEM[1759] + MEM[17462];
assign MEM[18192] = MEM[1762] + MEM[7456];
assign MEM[18193] = MEM[1763] + MEM[12410];
assign MEM[18194] = MEM[1764] + MEM[7391];
assign MEM[18195] = MEM[1767] + MEM[9291];
assign MEM[18196] = MEM[1771] + MEM[1851];
assign MEM[18197] = MEM[1772] + MEM[3876];
assign MEM[18198] = MEM[1773] + MEM[8566];
assign MEM[18199] = MEM[1774] + MEM[13652];
assign MEM[18200] = MEM[1775] + MEM[13546];
assign MEM[18201] = MEM[1780] + MEM[13001];
assign MEM[18202] = MEM[1781] + MEM[7994];
assign MEM[18203] = MEM[1782] + MEM[12056];
assign MEM[18204] = MEM[1790] + MEM[13133];
assign MEM[18205] = MEM[1791] + MEM[5111];
assign MEM[18206] = MEM[1803] + MEM[13026];
assign MEM[18207] = MEM[1804] + MEM[14961];
assign MEM[18208] = MEM[1805] + MEM[7727];
assign MEM[18209] = MEM[1806] + MEM[3949];
assign MEM[18210] = MEM[1811] + MEM[7577];
assign MEM[18211] = MEM[1813] + MEM[14230];
assign MEM[18212] = MEM[1814] + MEM[9524];
assign MEM[18213] = MEM[1815] + MEM[5738];
assign MEM[18214] = MEM[1818] + MEM[9346];
assign MEM[18215] = MEM[1820] + MEM[6111];
assign MEM[18216] = MEM[1821] + MEM[8363];
assign MEM[18217] = MEM[1822] + MEM[12918];
assign MEM[18218] = MEM[1826] + MEM[11150];
assign MEM[18219] = MEM[1827] + MEM[3245];
assign MEM[18220] = MEM[1828] + MEM[6171];
assign MEM[18221] = MEM[1829] + MEM[13597];
assign MEM[18222] = MEM[1830] + MEM[4858];
assign MEM[18223] = MEM[1835] + MEM[6707];
assign MEM[18224] = MEM[1836] + MEM[2908];
assign MEM[18225] = MEM[1837] + MEM[14226];
assign MEM[18226] = MEM[1838] + MEM[3916];
assign MEM[18227] = MEM[1843] + MEM[4951];
assign MEM[18228] = MEM[1844] + MEM[13202];
assign MEM[18229] = MEM[1845] + MEM[2447];
assign MEM[18230] = MEM[1846] + MEM[7366];
assign MEM[18231] = MEM[1852] + MEM[11141];
assign MEM[18232] = MEM[1854] + MEM[7484];
assign MEM[18233] = MEM[1859] + MEM[4386];
assign MEM[18234] = MEM[1860] + MEM[6276];
assign MEM[18235] = MEM[1861] + MEM[5813];
assign MEM[18236] = MEM[1867] + MEM[13050];
assign MEM[18237] = MEM[1868] + MEM[2527];
assign MEM[18238] = MEM[1869] + MEM[2238];
assign MEM[18239] = MEM[1875] + MEM[14999];
assign MEM[18240] = MEM[1877] + MEM[12267];
assign MEM[18241] = MEM[1878] + MEM[4271];
assign MEM[18242] = MEM[1879] + MEM[13627];
assign MEM[18243] = MEM[1882] + MEM[5635];
assign MEM[18244] = MEM[1883] + MEM[4911];
assign MEM[18245] = MEM[1884] + MEM[5119];
assign MEM[18246] = MEM[1885] + MEM[7909];
assign MEM[18247] = MEM[1886] + MEM[1927];
assign MEM[18248] = MEM[1887] + MEM[10765];
assign MEM[18249] = MEM[1891] + MEM[9029];
assign MEM[18250] = MEM[1893] + MEM[3076];
assign MEM[18251] = MEM[1895] + MEM[12342];
assign MEM[18252] = MEM[1899] + MEM[14968];
assign MEM[18253] = MEM[1901] + MEM[5356];
assign MEM[18254] = MEM[1903] + MEM[6586];
assign MEM[18255] = MEM[1907] + MEM[7647];
assign MEM[18256] = MEM[1909] + MEM[2100];
assign MEM[18257] = MEM[1910] + MEM[7768];
assign MEM[18258] = MEM[1914] + MEM[3149];
assign MEM[18259] = MEM[1915] + MEM[7285];
assign MEM[18260] = MEM[1917] + MEM[7304];
assign MEM[18261] = MEM[1918] + MEM[3890];
assign MEM[18262] = MEM[1922] + MEM[11056];
assign MEM[18263] = MEM[1925] + MEM[13307];
assign MEM[18264] = MEM[1932] + MEM[12428];
assign MEM[18265] = MEM[1933] + MEM[3671];
assign MEM[18266] = MEM[1935] + MEM[2294];
assign MEM[18267] = MEM[1938] + MEM[12108];
assign MEM[18268] = MEM[1939] + MEM[12541];
assign MEM[18269] = MEM[1949] + MEM[5894];
assign MEM[18270] = MEM[1950] + MEM[12249];
assign MEM[18271] = MEM[1951] + MEM[10947];
assign MEM[18272] = MEM[1954] + MEM[4542];
assign MEM[18273] = MEM[1955] + MEM[6718];
assign MEM[18274] = MEM[1956] + MEM[12150];
assign MEM[18275] = MEM[1957] + MEM[4126];
assign MEM[18276] = MEM[1962] + MEM[2509];
assign MEM[18277] = MEM[1965] + MEM[14683];
assign MEM[18278] = MEM[1966] + MEM[7152];
assign MEM[18279] = MEM[1967] + MEM[3732];
assign MEM[18280] = MEM[1970] + MEM[12222];
assign MEM[18281] = MEM[1971] + MEM[3101];
assign MEM[18282] = MEM[1975] + MEM[3027];
assign MEM[18283] = MEM[1978] + MEM[9657];
assign MEM[18284] = MEM[1979] + MEM[8000];
assign MEM[18285] = MEM[1980] + MEM[3038];
assign MEM[18286] = MEM[1981] + MEM[9006];
assign MEM[18287] = MEM[1982] + MEM[12432];
assign MEM[18288] = MEM[1983] + MEM[8088];
assign MEM[18289] = MEM[1984] + MEM[4716];
assign MEM[18290] = MEM[1986] + MEM[12091];
assign MEM[18291] = MEM[1987] + MEM[5087];
assign MEM[18292] = MEM[1989] + MEM[9707];
assign MEM[18293] = MEM[1990] + MEM[12584];
assign MEM[18294] = MEM[1991] + MEM[3781];
assign MEM[18295] = MEM[1995] + MEM[4615];
assign MEM[18296] = MEM[1997] + MEM[10760];
assign MEM[18297] = MEM[1998] + MEM[12784];
assign MEM[18298] = MEM[2002] + MEM[3725];
assign MEM[18299] = MEM[2003] + MEM[4091];
assign MEM[18300] = MEM[2004] + MEM[7738];
assign MEM[18301] = MEM[2005] + MEM[3485];
assign MEM[18302] = MEM[2011] + MEM[13313];
assign MEM[18303] = MEM[2013] + MEM[10466];
assign MEM[18304] = MEM[2014] + MEM[4077];
assign MEM[18305] = MEM[2023] + MEM[4111];
assign MEM[18306] = MEM[2031] + MEM[13054];
assign MEM[18307] = MEM[2034] + MEM[3693];
assign MEM[18308] = MEM[2035] + MEM[2684];
assign MEM[18309] = MEM[2036] + MEM[10589];
assign MEM[18310] = MEM[2037] + MEM[4524];
assign MEM[18311] = MEM[2039] + MEM[17285];
assign MEM[18312] = MEM[2042] + MEM[13708];
assign MEM[18313] = MEM[2043] + MEM[10019];
assign MEM[18314] = MEM[2045] + MEM[14913];
assign MEM[18315] = MEM[2046] + MEM[14852];
assign MEM[18316] = MEM[2050] + MEM[9799];
assign MEM[18317] = MEM[2052] + MEM[10746];
assign MEM[18318] = MEM[2053] + MEM[6422];
assign MEM[18319] = MEM[2054] + MEM[16540];
assign MEM[18320] = MEM[2058] + MEM[2146];
assign MEM[18321] = MEM[2060] + MEM[15221];
assign MEM[18322] = MEM[2061] + MEM[2211];
assign MEM[18323] = MEM[2062] + MEM[7502];
assign MEM[18324] = MEM[2070] + MEM[6464];
assign MEM[18325] = MEM[2075] + MEM[5660];
assign MEM[18326] = MEM[2077] + MEM[15319];
assign MEM[18327] = MEM[2082] + MEM[2443];
assign MEM[18328] = MEM[2083] + MEM[4006];
assign MEM[18329] = MEM[2086] + MEM[6037];
assign MEM[18330] = MEM[2087] + MEM[4302];
assign MEM[18331] = MEM[2090] + MEM[8020];
assign MEM[18332] = MEM[2091] + MEM[4509];
assign MEM[18333] = MEM[2093] + MEM[14651];
assign MEM[18334] = MEM[2095] + MEM[9077];
assign MEM[18335] = MEM[2101] + MEM[7332];
assign MEM[18336] = MEM[2102] + MEM[5839];
assign MEM[18337] = MEM[2109] + MEM[8090];
assign MEM[18338] = MEM[2116] + MEM[4058];
assign MEM[18339] = MEM[2124] + MEM[6904];
assign MEM[18340] = MEM[2125] + MEM[2140];
assign MEM[18341] = MEM[2126] + MEM[3476];
assign MEM[18342] = MEM[2130] + MEM[8295];
assign MEM[18343] = MEM[2133] + MEM[6442];
assign MEM[18344] = MEM[2135] + MEM[16973];
assign MEM[18345] = MEM[2138] + MEM[9350];
assign MEM[18346] = MEM[2139] + MEM[3877];
assign MEM[18347] = MEM[2147] + MEM[4334];
assign MEM[18348] = MEM[2148] + MEM[6343];
assign MEM[18349] = MEM[2154] + MEM[9547];
assign MEM[18350] = MEM[2156] + MEM[12294];
assign MEM[18351] = MEM[2157] + MEM[5021];
assign MEM[18352] = MEM[2159] + MEM[6130];
assign MEM[18353] = MEM[2163] + MEM[8384];
assign MEM[18354] = MEM[2165] + MEM[4287];
assign MEM[18355] = MEM[2167] + MEM[5295];
assign MEM[18356] = MEM[2170] + MEM[8470];
assign MEM[18357] = MEM[2172] + MEM[6905];
assign MEM[18358] = MEM[2173] + MEM[13266];
assign MEM[18359] = MEM[2175] + MEM[3292];
assign MEM[18360] = MEM[2178] + MEM[4090];
assign MEM[18361] = MEM[2179] + MEM[8008];
assign MEM[18362] = MEM[2181] + MEM[6635];
assign MEM[18363] = MEM[2183] + MEM[11343];
assign MEM[18364] = MEM[2186] + MEM[9187];
assign MEM[18365] = MEM[2189] + MEM[12484];
assign MEM[18366] = MEM[2194] + MEM[2303];
assign MEM[18367] = MEM[2195] + MEM[3607];
assign MEM[18368] = MEM[2198] + MEM[13912];
assign MEM[18369] = MEM[2199] + MEM[3572];
assign MEM[18370] = MEM[2203] + MEM[9873];
assign MEM[18371] = MEM[2204] + MEM[3202];
assign MEM[18372] = MEM[2207] + MEM[10742];
assign MEM[18373] = MEM[2210] + MEM[7615];
assign MEM[18374] = MEM[2212] + MEM[12936];
assign MEM[18375] = MEM[2214] + MEM[2957];
assign MEM[18376] = MEM[2215] + MEM[8043];
assign MEM[18377] = MEM[2226] + MEM[2679];
assign MEM[18378] = MEM[2230] + MEM[10507];
assign MEM[18379] = MEM[2231] + MEM[3756];
assign MEM[18380] = MEM[2235] + MEM[14193];
assign MEM[18381] = MEM[2237] + MEM[2635];
assign MEM[18382] = MEM[2239] + MEM[7595];
assign MEM[18383] = MEM[2246] + MEM[7324];
assign MEM[18384] = MEM[2247] + MEM[12593];
assign MEM[18385] = MEM[2252] + MEM[11215];
assign MEM[18386] = MEM[2255] + MEM[3116];
assign MEM[18387] = MEM[2260] + MEM[5702];
assign MEM[18388] = MEM[2261] + MEM[3534];
assign MEM[18389] = MEM[2267] + MEM[4262];
assign MEM[18390] = MEM[2268] + MEM[2673];
assign MEM[18391] = MEM[2270] + MEM[10828];
assign MEM[18392] = MEM[2271] + MEM[3516];
assign MEM[18393] = MEM[2285] + MEM[11136];
assign MEM[18394] = MEM[2286] + MEM[5661];
assign MEM[18395] = MEM[2287] + MEM[17363];
assign MEM[18396] = MEM[2292] + MEM[12113];
assign MEM[18397] = MEM[2298] + MEM[8603];
assign MEM[18398] = MEM[2299] + MEM[5140];
assign MEM[18399] = MEM[2300] + MEM[12524];
assign MEM[18400] = MEM[2308] + MEM[6969];
assign MEM[18401] = MEM[2310] + MEM[13803];
assign MEM[18402] = MEM[2314] + MEM[15073];
assign MEM[18403] = MEM[2315] + MEM[10287];
assign MEM[18404] = MEM[2317] + MEM[7130];
assign MEM[18405] = MEM[2318] + MEM[4198];
assign MEM[18406] = MEM[2319] + MEM[7579];
assign MEM[18407] = MEM[2324] + MEM[12650];
assign MEM[18408] = MEM[2330] + MEM[9363];
assign MEM[18409] = MEM[2331] + MEM[12717];
assign MEM[18410] = MEM[2334] + MEM[14254];
assign MEM[18411] = MEM[2338] + MEM[8249];
assign MEM[18412] = MEM[2341] + MEM[8838];
assign MEM[18413] = MEM[2342] + MEM[13109];
assign MEM[18414] = MEM[2343] + MEM[6881];
assign MEM[18415] = MEM[2347] + MEM[13408];
assign MEM[18416] = MEM[2348] + MEM[11312];
assign MEM[18417] = MEM[2349] + MEM[10856];
assign MEM[18418] = MEM[2354] + MEM[12465];
assign MEM[18419] = MEM[2355] + MEM[3034];
assign MEM[18420] = MEM[2356] + MEM[7594];
assign MEM[18421] = MEM[2358] + MEM[3374];
assign MEM[18422] = MEM[2367] + MEM[8386];
assign MEM[18423] = MEM[2371] + MEM[13148];
assign MEM[18424] = MEM[2373] + MEM[10983];
assign MEM[18425] = MEM[2374] + MEM[14339];
assign MEM[18426] = MEM[2375] + MEM[2839];
assign MEM[18427] = MEM[2379] + MEM[9357];
assign MEM[18428] = MEM[2381] + MEM[13783];
assign MEM[18429] = MEM[2382] + MEM[10775];
assign MEM[18430] = MEM[2383] + MEM[4210];
assign MEM[18431] = MEM[2386] + MEM[4421];
assign MEM[18432] = MEM[2387] + MEM[2867];
assign MEM[18433] = MEM[2389] + MEM[13306];
assign MEM[18434] = MEM[2391] + MEM[3127];
assign MEM[18435] = MEM[2394] + MEM[2831];
assign MEM[18436] = MEM[2396] + MEM[10115];
assign MEM[18437] = MEM[2405] + MEM[3914];
assign MEM[18438] = MEM[2411] + MEM[8958];
assign MEM[18439] = MEM[2413] + MEM[4580];
assign MEM[18440] = MEM[2415] + MEM[6220];
assign MEM[18441] = MEM[2418] + MEM[10743];
assign MEM[18442] = MEM[2419] + MEM[12333];
assign MEM[18443] = MEM[2420] + MEM[10643];
assign MEM[18444] = MEM[2422] + MEM[2543];
assign MEM[18445] = MEM[2426] + MEM[13690];
assign MEM[18446] = MEM[2427] + MEM[12450];
assign MEM[18447] = MEM[2429] + MEM[9182];
assign MEM[18448] = MEM[2430] + MEM[6262];
assign MEM[18449] = MEM[2431] + MEM[4202];
assign MEM[18450] = MEM[2434] + MEM[6124];
assign MEM[18451] = MEM[2435] + MEM[5524];
assign MEM[18452] = MEM[2437] + MEM[13870];
assign MEM[18453] = MEM[2438] + MEM[12126];
assign MEM[18454] = MEM[2442] + MEM[4511];
assign MEM[18455] = MEM[2444] + MEM[3959];
assign MEM[18456] = MEM[2450] + MEM[15398];
assign MEM[18457] = MEM[2451] + MEM[11090];
assign MEM[18458] = MEM[2452] + MEM[11662];
assign MEM[18459] = MEM[2453] + MEM[3652];
assign MEM[18460] = MEM[2462] + MEM[11210];
assign MEM[18461] = MEM[2463] + MEM[8906];
assign MEM[18462] = MEM[2468] + MEM[5067];
assign MEM[18463] = MEM[2469] + MEM[6570];
assign MEM[18464] = MEM[2471] + MEM[4172];
assign MEM[18465] = MEM[2475] + MEM[2988];
assign MEM[18466] = MEM[2477] + MEM[8762];
assign MEM[18467] = MEM[2478] + MEM[10909];
assign MEM[18468] = MEM[2479] + MEM[6139];
assign MEM[18469] = MEM[2486] + MEM[14264];
assign MEM[18470] = MEM[2487] + MEM[15368];
assign MEM[18471] = MEM[2490] + MEM[11976];
assign MEM[18472] = MEM[2500] + MEM[6964];
assign MEM[18473] = MEM[2501] + MEM[7754];
assign MEM[18474] = MEM[2502] + MEM[12765];
assign MEM[18475] = MEM[2508] + MEM[3884];
assign MEM[18476] = MEM[2510] + MEM[6923];
assign MEM[18477] = MEM[2511] + MEM[10024];
assign MEM[18478] = MEM[2514] + MEM[4835];
assign MEM[18479] = MEM[2516] + MEM[3308];
assign MEM[18480] = MEM[2517] + MEM[2943];
assign MEM[18481] = MEM[2522] + MEM[5899];
assign MEM[18482] = MEM[2524] + MEM[8769];
assign MEM[18483] = MEM[2526] + MEM[10943];
assign MEM[18484] = MEM[2530] + MEM[12227];
assign MEM[18485] = MEM[2531] + MEM[14219];
assign MEM[18486] = MEM[2532] + MEM[5591];
assign MEM[18487] = MEM[2533] + MEM[4772];
assign MEM[18488] = MEM[2538] + MEM[11954];
assign MEM[18489] = MEM[2539] + MEM[8564];
assign MEM[18490] = MEM[2540] + MEM[5487];
assign MEM[18491] = MEM[2541] + MEM[6661];
assign MEM[18492] = MEM[2548] + MEM[4730];
assign MEM[18493] = MEM[2558] + MEM[8671];
assign MEM[18494] = MEM[2562] + MEM[7120];
assign MEM[18495] = MEM[2564] + MEM[11012];
assign MEM[18496] = MEM[2567] + MEM[7877];
assign MEM[18497] = MEM[2570] + MEM[5102];
assign MEM[18498] = MEM[2571] + MEM[6125];
assign MEM[18499] = MEM[2573] + MEM[4614];
assign MEM[18500] = MEM[2574] + MEM[3446];
assign MEM[18501] = MEM[2581] + MEM[3066];
assign MEM[18502] = MEM[2586] + MEM[9343];
assign MEM[18503] = MEM[2588] + MEM[5735];
assign MEM[18504] = MEM[2594] + MEM[5420];
assign MEM[18505] = MEM[2595] + MEM[4340];
assign MEM[18506] = MEM[2598] + MEM[7517];
assign MEM[18507] = MEM[2599] + MEM[7438];
assign MEM[18508] = MEM[2602] + MEM[12684];
assign MEM[18509] = MEM[2604] + MEM[9733];
assign MEM[18510] = MEM[2605] + MEM[11310];
assign MEM[18511] = MEM[2606] + MEM[12425];
assign MEM[18512] = MEM[2607] + MEM[8439];
assign MEM[18513] = MEM[2610] + MEM[13170];
assign MEM[18514] = MEM[2611] + MEM[9311];
assign MEM[18515] = MEM[2613] + MEM[4479];
assign MEM[18516] = MEM[2615] + MEM[2623];
assign MEM[18517] = MEM[2618] + MEM[10918];
assign MEM[18518] = MEM[2620] + MEM[9487];
assign MEM[18519] = MEM[2622] + MEM[13949];
assign MEM[18520] = MEM[2630] + MEM[7247];
assign MEM[18521] = MEM[2636] + MEM[2818];
assign MEM[18522] = MEM[2638] + MEM[8643];
assign MEM[18523] = MEM[2639] + MEM[5870];
assign MEM[18524] = MEM[2643] + MEM[9244];
assign MEM[18525] = MEM[2645] + MEM[12156];
assign MEM[18526] = MEM[2647] + MEM[3206];
assign MEM[18527] = MEM[2650] + MEM[3924];
assign MEM[18528] = MEM[2655] + MEM[4796];
assign MEM[18529] = MEM[2657] + MEM[5690];
assign MEM[18530] = MEM[2658] + MEM[4285];
assign MEM[18531] = MEM[2661] + MEM[5634];
assign MEM[18532] = MEM[2662] + MEM[5530];
assign MEM[18533] = MEM[2663] + MEM[13644];
assign MEM[18534] = MEM[2665] + MEM[12413];
assign MEM[18535] = MEM[2668] + MEM[12337];
assign MEM[18536] = MEM[2669] + MEM[12805];
assign MEM[18537] = MEM[2671] + MEM[6837];
assign MEM[18538] = MEM[2672] + MEM[4332];
assign MEM[18539] = MEM[2674] + MEM[4469];
assign MEM[18540] = MEM[2676] + MEM[11374];
assign MEM[18541] = MEM[2677] + MEM[10230];
assign MEM[18542] = MEM[2685] + MEM[9401];
assign MEM[18543] = MEM[2687] + MEM[9462];
assign MEM[18544] = MEM[2692] + MEM[10791];
assign MEM[18545] = MEM[2693] + MEM[5782];
assign MEM[18546] = MEM[2694] + MEM[12576];
assign MEM[18547] = MEM[2699] + MEM[3660];
assign MEM[18548] = MEM[2700] + MEM[14514];
assign MEM[18549] = MEM[2702] + MEM[2789];
assign MEM[18550] = MEM[2703] + MEM[9841];
assign MEM[18551] = MEM[2706] + MEM[7656];
assign MEM[18552] = MEM[2707] + MEM[12426];
assign MEM[18553] = MEM[2708] + MEM[10675];
assign MEM[18554] = MEM[2715] + MEM[9608];
assign MEM[18555] = MEM[2716] + MEM[10916];
assign MEM[18556] = MEM[2724] + MEM[8461];
assign MEM[18557] = MEM[2727] + MEM[11254];
assign MEM[18558] = MEM[2730] + MEM[5196];
assign MEM[18559] = MEM[2734] + MEM[8204];
assign MEM[18560] = MEM[2735] + MEM[5301];
assign MEM[18561] = MEM[2740] + MEM[10621];
assign MEM[18562] = MEM[2741] + MEM[2802];
assign MEM[18563] = MEM[2742] + MEM[5316];
assign MEM[18564] = MEM[2744] + MEM[6821];
assign MEM[18565] = MEM[2750] + MEM[9034];
assign MEM[18566] = MEM[2751] + MEM[8998];
assign MEM[18567] = MEM[2754] + MEM[4683];
assign MEM[18568] = MEM[2755] + MEM[10800];
assign MEM[18569] = MEM[2756] + MEM[4765];
assign MEM[18570] = MEM[2757] + MEM[3874];
assign MEM[18571] = MEM[2758] + MEM[9651];
assign MEM[18572] = MEM[2759] + MEM[5313];
assign MEM[18573] = MEM[2762] + MEM[15752];
assign MEM[18574] = MEM[2764] + MEM[12804];
assign MEM[18575] = MEM[2765] + MEM[8182];
assign MEM[18576] = MEM[2766] + MEM[12578];
assign MEM[18577] = MEM[2770] + MEM[2946];
assign MEM[18578] = MEM[2774] + MEM[4014];
assign MEM[18579] = MEM[2775] + MEM[6976];
assign MEM[18580] = MEM[2779] + MEM[4692];
assign MEM[18581] = MEM[2781] + MEM[8942];
assign MEM[18582] = MEM[2783] + MEM[3052];
assign MEM[18583] = MEM[2786] + MEM[6823];
assign MEM[18584] = MEM[2787] + MEM[11352];
assign MEM[18585] = MEM[2788] + MEM[12099];
assign MEM[18586] = MEM[2791] + MEM[13790];
assign MEM[18587] = MEM[2794] + MEM[11402];
assign MEM[18588] = MEM[2795] + MEM[6181];
assign MEM[18589] = MEM[2796] + MEM[10477];
assign MEM[18590] = MEM[2797] + MEM[8734];
assign MEM[18591] = MEM[2803] + MEM[4406];
assign MEM[18592] = MEM[2805] + MEM[15405];
assign MEM[18593] = MEM[2806] + MEM[7519];
assign MEM[18594] = MEM[2807] + MEM[11637];
assign MEM[18595] = MEM[2810] + MEM[7950];
assign MEM[18596] = MEM[2813] + MEM[15558];
assign MEM[18597] = MEM[2814] + MEM[6571];
assign MEM[18598] = MEM[2819] + MEM[5365];
assign MEM[18599] = MEM[2821] + MEM[5998];
assign MEM[18600] = MEM[2822] + MEM[12527];
assign MEM[18601] = MEM[2827] + MEM[3909];
assign MEM[18602] = MEM[2828] + MEM[3647];
assign MEM[18603] = MEM[2829] + MEM[12953];
assign MEM[18604] = MEM[2834] + MEM[12860];
assign MEM[18605] = MEM[2836] + MEM[12574];
assign MEM[18606] = MEM[2837] + MEM[7450];
assign MEM[18607] = MEM[2838] + MEM[13501];
assign MEM[18608] = MEM[2842] + MEM[12280];
assign MEM[18609] = MEM[2844] + MEM[3503];
assign MEM[18610] = MEM[2845] + MEM[6618];
assign MEM[18611] = MEM[2851] + MEM[7440];
assign MEM[18612] = MEM[2852] + MEM[8458];
assign MEM[18613] = MEM[2853] + MEM[12288];
assign MEM[18614] = MEM[2854] + MEM[13117];
assign MEM[18615] = MEM[2855] + MEM[12767];
assign MEM[18616] = MEM[2859] + MEM[12327];
assign MEM[18617] = MEM[2860] + MEM[6810];
assign MEM[18618] = MEM[2861] + MEM[4165];
assign MEM[18619] = MEM[2862] + MEM[13639];
assign MEM[18620] = MEM[2868] + MEM[6660];
assign MEM[18621] = MEM[2870] + MEM[3119];
assign MEM[18622] = MEM[2871] + MEM[2987];
assign MEM[18623] = MEM[2872] + MEM[3096];
assign MEM[18624] = MEM[2874] + MEM[11801];
assign MEM[18625] = MEM[2875] + MEM[3059];
assign MEM[18626] = MEM[2876] + MEM[10842];
assign MEM[18627] = MEM[2877] + MEM[7916];
assign MEM[18628] = MEM[2880] + MEM[4839];
assign MEM[18629] = MEM[2883] + MEM[8717];
assign MEM[18630] = MEM[2884] + MEM[3999];
assign MEM[18631] = MEM[2885] + MEM[5302];
assign MEM[18632] = MEM[2886] + MEM[4322];
assign MEM[18633] = MEM[2890] + MEM[11646];
assign MEM[18634] = MEM[2891] + MEM[12493];
assign MEM[18635] = MEM[2894] + MEM[3970];
assign MEM[18636] = MEM[2899] + MEM[4373];
assign MEM[18637] = MEM[2900] + MEM[11069];
assign MEM[18638] = MEM[2901] + MEM[9552];
assign MEM[18639] = MEM[2902] + MEM[6846];
assign MEM[18640] = MEM[2911] + MEM[6410];
assign MEM[18641] = MEM[2917] + MEM[12414];
assign MEM[18642] = MEM[2918] + MEM[13856];
assign MEM[18643] = MEM[2919] + MEM[7180];
assign MEM[18644] = MEM[2924] + MEM[10282];
assign MEM[18645] = MEM[2925] + MEM[6888];
assign MEM[18646] = MEM[2926] + MEM[8060];
assign MEM[18647] = MEM[2927] + MEM[4207];
assign MEM[18648] = MEM[2931] + MEM[7766];
assign MEM[18649] = MEM[2933] + MEM[4653];
assign MEM[18650] = MEM[2935] + MEM[3915];
assign MEM[18651] = MEM[2938] + MEM[7212];
assign MEM[18652] = MEM[2940] + MEM[8646];
assign MEM[18653] = MEM[2941] + MEM[3863];
assign MEM[18654] = MEM[2942] + MEM[13476];
assign MEM[18655] = MEM[2947] + MEM[12401];
assign MEM[18656] = MEM[2949] + MEM[3035];
assign MEM[18657] = MEM[2959] + MEM[3124];
assign MEM[18658] = MEM[2964] + MEM[12171];
assign MEM[18659] = MEM[2965] + MEM[8992];
assign MEM[18660] = MEM[2966] + MEM[6617];
assign MEM[18661] = MEM[2967] + MEM[9033];
assign MEM[18662] = MEM[2970] + MEM[3983];
assign MEM[18663] = MEM[2972] + MEM[13229];
assign MEM[18664] = MEM[2973] + MEM[3663];
assign MEM[18665] = MEM[2975] + MEM[5202];
assign MEM[18666] = MEM[2979] + MEM[11253];
assign MEM[18667] = MEM[2986] + MEM[3090];
assign MEM[18668] = MEM[2994] + MEM[13550];
assign MEM[18669] = MEM[2995] + MEM[5562];
assign MEM[18670] = MEM[2998] + MEM[7423];
assign MEM[18671] = MEM[3006] + MEM[6127];
assign MEM[18672] = MEM[3007] + MEM[8187];
assign MEM[18673] = MEM[3011] + MEM[6686];
assign MEM[18674] = MEM[3012] + MEM[13669];
assign MEM[18675] = MEM[3013] + MEM[3383];
assign MEM[18676] = MEM[3015] + MEM[12626];
assign MEM[18677] = MEM[3019] + MEM[5910];
assign MEM[18678] = MEM[3020] + MEM[3479];
assign MEM[18679] = MEM[3021] + MEM[10611];
assign MEM[18680] = MEM[3022] + MEM[5860];
assign MEM[18681] = MEM[3028] + MEM[8578];
assign MEM[18682] = MEM[3031] + MEM[12455];
assign MEM[18683] = MEM[3036] + MEM[4118];
assign MEM[18684] = MEM[3042] + MEM[4451];
assign MEM[18685] = MEM[3043] + MEM[3427];
assign MEM[18686] = MEM[3044] + MEM[3114];
assign MEM[18687] = MEM[3051] + MEM[10006];
assign MEM[18688] = MEM[3054] + MEM[12031];
assign MEM[18689] = MEM[3060] + MEM[13943];
assign MEM[18690] = MEM[3061] + MEM[5374];
assign MEM[18691] = MEM[3062] + MEM[12147];
assign MEM[18692] = MEM[3067] + MEM[13660];
assign MEM[18693] = MEM[3068] + MEM[14829];
assign MEM[18694] = MEM[3071] + MEM[6961];
assign MEM[18695] = MEM[3074] + MEM[7465];
assign MEM[18696] = MEM[3075] + MEM[7073];
assign MEM[18697] = MEM[3077] + MEM[12852];
assign MEM[18698] = MEM[3078] + MEM[11647];
assign MEM[18699] = MEM[3083] + MEM[5973];
assign MEM[18700] = MEM[3085] + MEM[11000];
assign MEM[18701] = MEM[3086] + MEM[14804];
assign MEM[18702] = MEM[3092] + MEM[9605];
assign MEM[18703] = MEM[3093] + MEM[14148];
assign MEM[18704] = MEM[3094] + MEM[5943];
assign MEM[18705] = MEM[3098] + MEM[7880];
assign MEM[18706] = MEM[3099] + MEM[13497];
assign MEM[18707] = MEM[3100] + MEM[5759];
assign MEM[18708] = MEM[3107] + MEM[13752];
assign MEM[18709] = MEM[3108] + MEM[12844];
assign MEM[18710] = MEM[3109] + MEM[12083];
assign MEM[18711] = MEM[3110] + MEM[3997];
assign MEM[18712] = MEM[3115] + MEM[9659];
assign MEM[18713] = MEM[3118] + MEM[5901];
assign MEM[18714] = MEM[3122] + MEM[3621];
assign MEM[18715] = MEM[3125] + MEM[4726];
assign MEM[18716] = MEM[3126] + MEM[7653];
assign MEM[18717] = MEM[3130] + MEM[14629];
assign MEM[18718] = MEM[3132] + MEM[7315];
assign MEM[18719] = MEM[3133] + MEM[17457];
assign MEM[18720] = MEM[3134] + MEM[4805];
assign MEM[18721] = MEM[3141] + MEM[5717];
assign MEM[18722] = MEM[3143] + MEM[4948];
assign MEM[18723] = MEM[3150] + MEM[3908];
assign MEM[18724] = MEM[3151] + MEM[9713];
assign MEM[18725] = MEM[3157] + MEM[4871];
assign MEM[18726] = MEM[3158] + MEM[9894];
assign MEM[18727] = MEM[3159] + MEM[4013];
assign MEM[18728] = MEM[3162] + MEM[13440];
assign MEM[18729] = MEM[3163] + MEM[3861];
assign MEM[18730] = MEM[3164] + MEM[8349];
assign MEM[18731] = MEM[3165] + MEM[5531];
assign MEM[18732] = MEM[3167] + MEM[3357];
assign MEM[18733] = MEM[3170] + MEM[7038];
assign MEM[18734] = MEM[3171] + MEM[10873];
assign MEM[18735] = MEM[3178] + MEM[7929];
assign MEM[18736] = MEM[3180] + MEM[5692];
assign MEM[18737] = MEM[3181] + MEM[12273];
assign MEM[18738] = MEM[3182] + MEM[10668];
assign MEM[18739] = MEM[3184] + MEM[13410];
assign MEM[18740] = MEM[3185] + MEM[10978];
assign MEM[18741] = MEM[3187] + MEM[13312];
assign MEM[18742] = MEM[3188] + MEM[12557];
assign MEM[18743] = MEM[3190] + MEM[14119];
assign MEM[18744] = MEM[3191] + MEM[11157];
assign MEM[18745] = MEM[3196] + MEM[8286];
assign MEM[18746] = MEM[3197] + MEM[11185];
assign MEM[18747] = MEM[3199] + MEM[6095];
assign MEM[18748] = MEM[3203] + MEM[7939];
assign MEM[18749] = MEM[3204] + MEM[7792];
assign MEM[18750] = MEM[3205] + MEM[3947];
assign MEM[18751] = MEM[3207] + MEM[11982];
assign MEM[18752] = MEM[3210] + MEM[4538];
assign MEM[18753] = MEM[3211] + MEM[15277];
assign MEM[18754] = MEM[3212] + MEM[13048];
assign MEM[18755] = MEM[3214] + MEM[6591];
assign MEM[18756] = MEM[3215] + MEM[3995];
assign MEM[18757] = MEM[3220] + MEM[12195];
assign MEM[18758] = MEM[3222] + MEM[7524];
assign MEM[18759] = MEM[3227] + MEM[9102];
assign MEM[18760] = MEM[3229] + MEM[5883];
assign MEM[18761] = MEM[3231] + MEM[3941];
assign MEM[18762] = MEM[3236] + MEM[5878];
assign MEM[18763] = MEM[3239] + MEM[3508];
assign MEM[18764] = MEM[3244] + MEM[4693];
assign MEM[18765] = MEM[3246] + MEM[6377];
assign MEM[18766] = MEM[3247] + MEM[9301];
assign MEM[18767] = MEM[3251] + MEM[13085];
assign MEM[18768] = MEM[3253] + MEM[7124];
assign MEM[18769] = MEM[3255] + MEM[13434];
assign MEM[18770] = MEM[3259] + MEM[5911];
assign MEM[18771] = MEM[3260] + MEM[4078];
assign MEM[18772] = MEM[3262] + MEM[10874];
assign MEM[18773] = MEM[3267] + MEM[3842];
assign MEM[18774] = MEM[3268] + MEM[4487];
assign MEM[18775] = MEM[3269] + MEM[15220];
assign MEM[18776] = MEM[3270] + MEM[6993];
assign MEM[18777] = MEM[3271] + MEM[12743];
assign MEM[18778] = MEM[3275] + MEM[12785];
assign MEM[18779] = MEM[3276] + MEM[10232];
assign MEM[18780] = MEM[3277] + MEM[9621];
assign MEM[18781] = MEM[3278] + MEM[10568];
assign MEM[18782] = MEM[3283] + MEM[4466];
assign MEM[18783] = MEM[3284] + MEM[5940];
assign MEM[18784] = MEM[3285] + MEM[13620];
assign MEM[18785] = MEM[3286] + MEM[8864];
assign MEM[18786] = MEM[3287] + MEM[10463];
assign MEM[18787] = MEM[3291] + MEM[11962];
assign MEM[18788] = MEM[3295] + MEM[3602];
assign MEM[18789] = MEM[3298] + MEM[12526];
assign MEM[18790] = MEM[3300] + MEM[3939];
assign MEM[18791] = MEM[3301] + MEM[12335];
assign MEM[18792] = MEM[3307] + MEM[7660];
assign MEM[18793] = MEM[3309] + MEM[12624];
assign MEM[18794] = MEM[3311] + MEM[12365];
assign MEM[18795] = MEM[3314] + MEM[4964];
assign MEM[18796] = MEM[3316] + MEM[10461];
assign MEM[18797] = MEM[3319] + MEM[12950];
assign MEM[18798] = MEM[3322] + MEM[11023];
assign MEM[18799] = MEM[3323] + MEM[5979];
assign MEM[18800] = MEM[3324] + MEM[11915];
assign MEM[18801] = MEM[3326] + MEM[16992];
assign MEM[18802] = MEM[3327] + MEM[4822];
assign MEM[18803] = MEM[3330] + MEM[6942];
assign MEM[18804] = MEM[3331] + MEM[8334];
assign MEM[18805] = MEM[3332] + MEM[7566];
assign MEM[18806] = MEM[3333] + MEM[10841];
assign MEM[18807] = MEM[3334] + MEM[8223];
assign MEM[18808] = MEM[3338] + MEM[4779];
assign MEM[18809] = MEM[3339] + MEM[5778];
assign MEM[18810] = MEM[3340] + MEM[3887];
assign MEM[18811] = MEM[3342] + MEM[5711];
assign MEM[18812] = MEM[3347] + MEM[12353];
assign MEM[18813] = MEM[3349] + MEM[9750];
assign MEM[18814] = MEM[3350] + MEM[3778];
assign MEM[18815] = MEM[3358] + MEM[16474];
assign MEM[18816] = MEM[3365] + MEM[8504];
assign MEM[18817] = MEM[3371] + MEM[8036];
assign MEM[18818] = MEM[3373] + MEM[14218];
assign MEM[18819] = MEM[3380] + MEM[7685];
assign MEM[18820] = MEM[3383] + MEM[9315];
assign MEM[18821] = MEM[3387] + MEM[4530];
assign MEM[18822] = MEM[3389] + MEM[7132];
assign MEM[18823] = MEM[3394] + MEM[3933];
assign MEM[18824] = MEM[3395] + MEM[9432];
assign MEM[18825] = MEM[3397] + MEM[4903];
assign MEM[18826] = MEM[3399] + MEM[4851];
assign MEM[18827] = MEM[3404] + MEM[11389];
assign MEM[18828] = MEM[3406] + MEM[5055];
assign MEM[18829] = MEM[3410] + MEM[15071];
assign MEM[18830] = MEM[3412] + MEM[6094];
assign MEM[18831] = MEM[3414] + MEM[8149];
assign MEM[18832] = MEM[3415] + MEM[13441];
assign MEM[18833] = MEM[3418] + MEM[12821];
assign MEM[18834] = MEM[3420] + MEM[11975];
assign MEM[18835] = MEM[3422] + MEM[7957];
assign MEM[18836] = MEM[3423] + MEM[13066];
assign MEM[18837] = MEM[3429] + MEM[6875];
assign MEM[18838] = MEM[3434] + MEM[5475];
assign MEM[18839] = MEM[3437] + MEM[11644];
assign MEM[18840] = MEM[3438] + MEM[8253];
assign MEM[18841] = MEM[3439] + MEM[7329];
assign MEM[18842] = MEM[3444] + MEM[4355];
assign MEM[18843] = MEM[3447] + MEM[7214];
assign MEM[18844] = MEM[3451] + MEM[4582];
assign MEM[18845] = MEM[3452] + MEM[7860];
assign MEM[18846] = MEM[3453] + MEM[8301];
assign MEM[18847] = MEM[3458] + MEM[7233];
assign MEM[18848] = MEM[3459] + MEM[9687];
assign MEM[18849] = MEM[3461] + MEM[4517];
assign MEM[18850] = MEM[3467] + MEM[4814];
assign MEM[18851] = MEM[3470] + MEM[10906];
assign MEM[18852] = MEM[3475] + MEM[11474];
assign MEM[18853] = MEM[3477] + MEM[10699];
assign MEM[18854] = MEM[3478] + MEM[4579];
assign MEM[18855] = MEM[3482] + MEM[8802];
assign MEM[18856] = MEM[3483] + MEM[14420];
assign MEM[18857] = MEM[3484] + MEM[12039];
assign MEM[18858] = MEM[3487] + MEM[4862];
assign MEM[18859] = MEM[3490] + MEM[13695];
assign MEM[18860] = MEM[3493] + MEM[13474];
assign MEM[18861] = MEM[3494] + MEM[11799];
assign MEM[18862] = MEM[3499] + MEM[12548];
assign MEM[18863] = MEM[3500] + MEM[5007];
assign MEM[18864] = MEM[3501] + MEM[12569];
assign MEM[18865] = MEM[3502] + MEM[11115];
assign MEM[18866] = MEM[3507] + MEM[7367];
assign MEM[18867] = MEM[3511] + MEM[15016];
assign MEM[18868] = MEM[3514] + MEM[12668];
assign MEM[18869] = MEM[3515] + MEM[3994];
assign MEM[18870] = MEM[3517] + MEM[6717];
assign MEM[18871] = MEM[3518] + MEM[5458];
assign MEM[18872] = MEM[3519] + MEM[5470];
assign MEM[18873] = MEM[3526] + MEM[5684];
assign MEM[18874] = MEM[3531] + MEM[13194];
assign MEM[18875] = MEM[3532] + MEM[14486];
assign MEM[18876] = MEM[3533] + MEM[7424];
assign MEM[18877] = MEM[3535] + MEM[12565];
assign MEM[18878] = MEM[3539] + MEM[6431];
assign MEM[18879] = MEM[3540] + MEM[9776];
assign MEM[18880] = MEM[3542] + MEM[5271];
assign MEM[18881] = MEM[3543] + MEM[15728];
assign MEM[18882] = MEM[3546] + MEM[12596];
assign MEM[18883] = MEM[3547] + MEM[8658];
assign MEM[18884] = MEM[3548] + MEM[4678];
assign MEM[18885] = MEM[3549] + MEM[3775];
assign MEM[18886] = MEM[3550] + MEM[5970];
assign MEM[18887] = MEM[3554] + MEM[9243];
assign MEM[18888] = MEM[3556] + MEM[12685];
assign MEM[18889] = MEM[3557] + MEM[15092];
assign MEM[18890] = MEM[3564] + MEM[13759];
assign MEM[18891] = MEM[3565] + MEM[12774];
assign MEM[18892] = MEM[3566] + MEM[7869];
assign MEM[18893] = MEM[3567] + MEM[13114];
assign MEM[18894] = MEM[3571] + MEM[6694];
assign MEM[18895] = MEM[3573] + MEM[8655];
assign MEM[18896] = MEM[3575] + MEM[11087];
assign MEM[18897] = MEM[3578] + MEM[8063];
assign MEM[18898] = MEM[3580] + MEM[10656];
assign MEM[18899] = MEM[3582] + MEM[12420];
assign MEM[18900] = MEM[3583] + MEM[4999];
assign MEM[18901] = MEM[3591] + MEM[15748];
assign MEM[18902] = MEM[3597] + MEM[11266];
assign MEM[18903] = MEM[3598] + MEM[6047];
assign MEM[18904] = MEM[3599] + MEM[4514];
assign MEM[18905] = MEM[3604] + MEM[3742];
assign MEM[18906] = MEM[3606] + MEM[13727];
assign MEM[18907] = MEM[3612] + MEM[12268];
assign MEM[18908] = MEM[3613] + MEM[8686];
assign MEM[18909] = MEM[3615] + MEM[13901];
assign MEM[18910] = MEM[3618] + MEM[12448];
assign MEM[18911] = MEM[3620] + MEM[4821];
assign MEM[18912] = MEM[3622] + MEM[8058];
assign MEM[18913] = MEM[3626] + MEM[3895];
assign MEM[18914] = MEM[3628] + MEM[8269];
assign MEM[18915] = MEM[3630] + MEM[5770];
assign MEM[18916] = MEM[3634] + MEM[12749];
assign MEM[18917] = MEM[3636] + MEM[6983];
assign MEM[18918] = MEM[3637] + MEM[5990];
assign MEM[18919] = MEM[3638] + MEM[11003];
assign MEM[18920] = MEM[3639] + MEM[10811];
assign MEM[18921] = MEM[3642] + MEM[4787];
assign MEM[18922] = MEM[3643] + MEM[7861];
assign MEM[18923] = MEM[3644] + MEM[12317];
assign MEM[18924] = MEM[3645] + MEM[5198];
assign MEM[18925] = MEM[3646] + MEM[5621];
assign MEM[18926] = MEM[3653] + MEM[8791];
assign MEM[18927] = MEM[3654] + MEM[7616];
assign MEM[18928] = MEM[3658] + MEM[7489];
assign MEM[18929] = MEM[3659] + MEM[7271];
assign MEM[18930] = MEM[3667] + MEM[5234];
assign MEM[18931] = MEM[3669] + MEM[4319];
assign MEM[18932] = MEM[3675] + MEM[13271];
assign MEM[18933] = MEM[3676] + MEM[14598];
assign MEM[18934] = MEM[3677] + MEM[7900];
assign MEM[18935] = MEM[3678] + MEM[7448];
assign MEM[18936] = MEM[3679] + MEM[10816];
assign MEM[18937] = MEM[3682] + MEM[4986];
assign MEM[18938] = MEM[3684] + MEM[13492];
assign MEM[18939] = MEM[3685] + MEM[8266];
assign MEM[18940] = MEM[3687] + MEM[15803];
assign MEM[18941] = MEM[3690] + MEM[7256];
assign MEM[18942] = MEM[3698] + MEM[10826];
assign MEM[18943] = MEM[3702] + MEM[9134];
assign MEM[18944] = MEM[3703] + MEM[8779];
assign MEM[18945] = MEM[3706] + MEM[15466];
assign MEM[18946] = MEM[3708] + MEM[4199];
assign MEM[18947] = MEM[3708] + MEM[9240];
assign MEM[18948] = MEM[3709] + MEM[10623];
assign MEM[18949] = MEM[3710] + MEM[7090];
assign MEM[18950] = MEM[3711] + MEM[9387];
assign MEM[18951] = MEM[3714] + MEM[9636];
assign MEM[18952] = MEM[3715] + MEM[6380];
assign MEM[18953] = MEM[3716] + MEM[3911];
assign MEM[18954] = MEM[3719] + MEM[8325];
assign MEM[18955] = MEM[3722] + MEM[7032];
assign MEM[18956] = MEM[3723] + MEM[9374];
assign MEM[18957] = MEM[3724] + MEM[14886];
assign MEM[18958] = MEM[3726] + MEM[14052];
assign MEM[18959] = MEM[3727] + MEM[12472];
assign MEM[18960] = MEM[3734] + MEM[5682];
assign MEM[18961] = MEM[3735] + MEM[4420];
assign MEM[18962] = MEM[3739] + MEM[10648];
assign MEM[18963] = MEM[3740] + MEM[4468];
assign MEM[18964] = MEM[3741] + MEM[3974];
assign MEM[18965] = MEM[3746] + MEM[4223];
assign MEM[18966] = MEM[3747] + MEM[5334];
assign MEM[18967] = MEM[3748] + MEM[7779];
assign MEM[18968] = MEM[3755] + MEM[8408];
assign MEM[18969] = MEM[3757] + MEM[7533];
assign MEM[18970] = MEM[3758] + MEM[7531];
assign MEM[18971] = MEM[3759] + MEM[13151];
assign MEM[18972] = MEM[3762] + MEM[9375];
assign MEM[18973] = MEM[3767] + MEM[12499];
assign MEM[18974] = MEM[3770] + MEM[12568];
assign MEM[18975] = MEM[3771] + MEM[4439];
assign MEM[18976] = MEM[3772] + MEM[5638];
assign MEM[18977] = MEM[3774] + MEM[10945];
assign MEM[18978] = MEM[3779] + MEM[14436];
assign MEM[18979] = MEM[3783] + MEM[7330];
assign MEM[18980] = MEM[3787] + MEM[7048];
assign MEM[18981] = MEM[3788] + MEM[6887];
assign MEM[18982] = MEM[3789] + MEM[7207];
assign MEM[18983] = MEM[3791] + MEM[8735];
assign MEM[18984] = MEM[3794] + MEM[5446];
assign MEM[18985] = MEM[3795] + MEM[9263];
assign MEM[18986] = MEM[3796] + MEM[13093];
assign MEM[18987] = MEM[3797] + MEM[3836];
assign MEM[18988] = MEM[3802] + MEM[13293];
assign MEM[18989] = MEM[3803] + MEM[12427];
assign MEM[18990] = MEM[3804] + MEM[6692];
assign MEM[18991] = MEM[3807] + MEM[11137];
assign MEM[18992] = MEM[3813] + MEM[5903];
assign MEM[18993] = MEM[3814] + MEM[5615];
assign MEM[18994] = MEM[3828] + MEM[4812];
assign MEM[18995] = MEM[3829] + MEM[5871];
assign MEM[18996] = MEM[3830] + MEM[14324];
assign MEM[18997] = MEM[3837] + MEM[9450];
assign MEM[18998] = MEM[3846] + MEM[11476];
assign MEM[18999] = MEM[3847] + MEM[4122];
assign MEM[19000] = MEM[3850] + MEM[7072];
assign MEM[19001] = MEM[3854] + MEM[11448];
assign MEM[19002] = MEM[3855] + MEM[5644];
assign MEM[19003] = MEM[3858] + MEM[12211];
assign MEM[19004] = MEM[3859] + MEM[5443];
assign MEM[19005] = MEM[3860] + MEM[5019];
assign MEM[19006] = MEM[3869] + MEM[11684];
assign MEM[19007] = MEM[3870] + MEM[12652];
assign MEM[19008] = MEM[3883] + MEM[4270];
assign MEM[19009] = MEM[3886] + MEM[7351];
assign MEM[19010] = MEM[3888] + MEM[3896];
assign MEM[19011] = MEM[3892] + MEM[11060];
assign MEM[19012] = MEM[3898] + MEM[11192];
assign MEM[19013] = MEM[3906] + MEM[10907];
assign MEM[19014] = MEM[3907] + MEM[8672];
assign MEM[19015] = MEM[3910] + MEM[7943];
assign MEM[19016] = MEM[3919] + MEM[5071];
assign MEM[19017] = MEM[3925] + MEM[9303];
assign MEM[19018] = MEM[3926] + MEM[5419];
assign MEM[19019] = MEM[3930] + MEM[13954];
assign MEM[19020] = MEM[3932] + MEM[12477];
assign MEM[19021] = MEM[3940] + MEM[4155];
assign MEM[19022] = MEM[3943] + MEM[5406];
assign MEM[19023] = MEM[3948] + MEM[6077];
assign MEM[19024] = MEM[3950] + MEM[16112];
assign MEM[19025] = MEM[3951] + MEM[9522];
assign MEM[19026] = MEM[3954] + MEM[14982];
assign MEM[19027] = MEM[3955] + MEM[4701];
assign MEM[19028] = MEM[3956] + MEM[7962];
assign MEM[19029] = MEM[3957] + MEM[5051];
assign MEM[19030] = MEM[3958] + MEM[12145];
assign MEM[19031] = MEM[3963] + MEM[6908];
assign MEM[19032] = MEM[3964] + MEM[12680];
assign MEM[19033] = MEM[3967] + MEM[4443];
assign MEM[19034] = MEM[3973] + MEM[8848];
assign MEM[19035] = MEM[3975] + MEM[7551];
assign MEM[19036] = MEM[3978] + MEM[7262];
assign MEM[19037] = MEM[3979] + MEM[9299];
assign MEM[19038] = MEM[3980] + MEM[4846];
assign MEM[19039] = MEM[3981] + MEM[6473];
assign MEM[19040] = MEM[3987] + MEM[7240];
assign MEM[19041] = MEM[3988] + MEM[11888];
assign MEM[19042] = MEM[3989] + MEM[4613];
assign MEM[19043] = MEM[3996] + MEM[4644];
assign MEM[19044] = MEM[3998] + MEM[13576];
assign MEM[19045] = MEM[4002] + MEM[10899];
assign MEM[19046] = MEM[4004] + MEM[13766];
assign MEM[19047] = MEM[4005] + MEM[9138];
assign MEM[19048] = MEM[4010] + MEM[9183];
assign MEM[19049] = MEM[4011] + MEM[4982];
assign MEM[19050] = MEM[4015] + MEM[7364];
assign MEM[19051] = MEM[4018] + MEM[10504];
assign MEM[19052] = MEM[4021] + MEM[9466];
assign MEM[19053] = MEM[4022] + MEM[5031];
assign MEM[19054] = MEM[4023] + MEM[4887];
assign MEM[19055] = MEM[4030] + MEM[8205];
assign MEM[19056] = MEM[4031] + MEM[11638];
assign MEM[19057] = MEM[4037] + MEM[8101];
assign MEM[19058] = MEM[4045] + MEM[6579];
assign MEM[19059] = MEM[4046] + MEM[4246];
assign MEM[19060] = MEM[4051] + MEM[9367];
assign MEM[19061] = MEM[4053] + MEM[11063];
assign MEM[19062] = MEM[4054] + MEM[11902];
assign MEM[19063] = MEM[4062] + MEM[8720];
assign MEM[19064] = MEM[4066] + MEM[10560];
assign MEM[19065] = MEM[4067] + MEM[6813];
assign MEM[19066] = MEM[4069] + MEM[10138];
assign MEM[19067] = MEM[4070] + MEM[10840];
assign MEM[19068] = MEM[4074] + MEM[11159];
assign MEM[19069] = MEM[4076] + MEM[6391];
assign MEM[19070] = MEM[4082] + MEM[8252];
assign MEM[19071] = MEM[4083] + MEM[4886];
assign MEM[19072] = MEM[4084] + MEM[12917];
assign MEM[19073] = MEM[4085] + MEM[11458];
assign MEM[19074] = MEM[4086] + MEM[10950];
assign MEM[19075] = MEM[4092] + MEM[6107];
assign MEM[19076] = MEM[4093] + MEM[11736];
assign MEM[19077] = MEM[4094] + MEM[8829];
assign MEM[19078] = MEM[4095] + MEM[7549];
assign MEM[19079] = MEM[4098] + MEM[4318];
assign MEM[19080] = MEM[4099] + MEM[7789];
assign MEM[19081] = MEM[4100] + MEM[8287];
assign MEM[19082] = MEM[4102] + MEM[9689];
assign MEM[19083] = MEM[4103] + MEM[4546];
assign MEM[19084] = MEM[4106] + MEM[7867];
assign MEM[19085] = MEM[4108] + MEM[6863];
assign MEM[19086] = MEM[4109] + MEM[6497];
assign MEM[19087] = MEM[4110] + MEM[9476];
assign MEM[19088] = MEM[4115] + MEM[7296];
assign MEM[19089] = MEM[4116] + MEM[12715];
assign MEM[19090] = MEM[4119] + MEM[12482];
assign MEM[19091] = MEM[4124] + MEM[15168];
assign MEM[19092] = MEM[4125] + MEM[12371];
assign MEM[19093] = MEM[4127] + MEM[12261];
assign MEM[19094] = MEM[4131] + MEM[6213];
assign MEM[19095] = MEM[4133] + MEM[12345];
assign MEM[19096] = MEM[4134] + MEM[13147];
assign MEM[19097] = MEM[4135] + MEM[4306];
assign MEM[19098] = MEM[4138] + MEM[11362];
assign MEM[19099] = MEM[4142] + MEM[7179];
assign MEM[19100] = MEM[4143] + MEM[4371];
assign MEM[19101] = MEM[4147] + MEM[7761];
assign MEM[19102] = MEM[4148] + MEM[14622];
assign MEM[19103] = MEM[4150] + MEM[6853];
assign MEM[19104] = MEM[4159] + MEM[5978];
assign MEM[19105] = MEM[4164] + MEM[4868];
assign MEM[19106] = MEM[4171] + MEM[11670];
assign MEM[19107] = MEM[4174] + MEM[6329];
assign MEM[19108] = MEM[4175] + MEM[10937];
assign MEM[19109] = MEM[4178] + MEM[15049];
assign MEM[19110] = MEM[4180] + MEM[17672];
assign MEM[19111] = MEM[4182] + MEM[7166];
assign MEM[19112] = MEM[4188] + MEM[12215];
assign MEM[19113] = MEM[4190] + MEM[14331];
assign MEM[19114] = MEM[4191] + MEM[12697];
assign MEM[19115] = MEM[4194] + MEM[7781];
assign MEM[19116] = MEM[4195] + MEM[10087];
assign MEM[19117] = MEM[4197] + MEM[13635];
assign MEM[19118] = MEM[4203] + MEM[8406];
assign MEM[19119] = MEM[4218] + MEM[12182];
assign MEM[19120] = MEM[4219] + MEM[11172];
assign MEM[19121] = MEM[4221] + MEM[17055];
assign MEM[19122] = MEM[4222] + MEM[12250];
assign MEM[19123] = MEM[4229] + MEM[5714];
assign MEM[19124] = MEM[4230] + MEM[14088];
assign MEM[19125] = MEM[4231] + MEM[6797];
assign MEM[19126] = MEM[4235] + MEM[4659];
assign MEM[19127] = MEM[4236] + MEM[7693];
assign MEM[19128] = MEM[4238] + MEM[8908];
assign MEM[19129] = MEM[4242] + MEM[7469];
assign MEM[19130] = MEM[4243] + MEM[10991];
assign MEM[19131] = MEM[4244] + MEM[7491];
assign MEM[19132] = MEM[4245] + MEM[12750];
assign MEM[19133] = MEM[4250] + MEM[11999];
assign MEM[19134] = MEM[4254] + MEM[13463];
assign MEM[19135] = MEM[4261] + MEM[8049];
assign MEM[19136] = MEM[4268] + MEM[5662];
assign MEM[19137] = MEM[4276] + MEM[12674];
assign MEM[19138] = MEM[4277] + MEM[8267];
assign MEM[19139] = MEM[4278] + MEM[13685];
assign MEM[19140] = MEM[4284] + MEM[7976];
assign MEM[19141] = MEM[4286] + MEM[13452];
assign MEM[19142] = MEM[4290] + MEM[10097];
assign MEM[19143] = MEM[4294] + MEM[11870];
assign MEM[19144] = MEM[4298] + MEM[5807];
assign MEM[19145] = MEM[4299] + MEM[7497];
assign MEM[19146] = MEM[4308] + MEM[11234];
assign MEM[19147] = MEM[4310] + MEM[5068];
assign MEM[19148] = MEM[4311] + MEM[6132];
assign MEM[19149] = MEM[4314] + MEM[12104];
assign MEM[19150] = MEM[4323] + MEM[5263];
assign MEM[19151] = MEM[4324] + MEM[4642];
assign MEM[19152] = MEM[4326] + MEM[8497];
assign MEM[19153] = MEM[4330] + MEM[11317];
assign MEM[19154] = MEM[4331] + MEM[10158];
assign MEM[19155] = MEM[4333] + MEM[7388];
assign MEM[19156] = MEM[4338] + MEM[14332];
assign MEM[19157] = MEM[4339] + MEM[10762];
assign MEM[19158] = MEM[4342] + MEM[10065];
assign MEM[19159] = MEM[4343] + MEM[4910];
assign MEM[19160] = MEM[4343] + MEM[13182];
assign MEM[19161] = MEM[4346] + MEM[14694];
assign MEM[19162] = MEM[4351] + MEM[8473];
assign MEM[19163] = MEM[4354] + MEM[8753];
assign MEM[19164] = MEM[4356] + MEM[9840];
assign MEM[19165] = MEM[4357] + MEM[9533];
assign MEM[19166] = MEM[4358] + MEM[4363];
assign MEM[19167] = MEM[4362] + MEM[16362];
assign MEM[19168] = MEM[4366] + MEM[9551];
assign MEM[19169] = MEM[4367] + MEM[6222];
assign MEM[19170] = MEM[4375] + MEM[16111];
assign MEM[19171] = MEM[4387] + MEM[7115];
assign MEM[19172] = MEM[4389] + MEM[12416];
assign MEM[19173] = MEM[4390] + MEM[12501];
assign MEM[19174] = MEM[4394] + MEM[6421];
assign MEM[19175] = MEM[4395] + MEM[12381];
assign MEM[19176] = MEM[4396] + MEM[9103];
assign MEM[19177] = MEM[4397] + MEM[15104];
assign MEM[19178] = MEM[4398] + MEM[9233];
assign MEM[19179] = MEM[4402] + MEM[6583];
assign MEM[19180] = MEM[4407] + MEM[11630];
assign MEM[19181] = MEM[4413] + MEM[4461];
assign MEM[19182] = MEM[4414] + MEM[4996];
assign MEM[19183] = MEM[4415] + MEM[6133];
assign MEM[19184] = MEM[4419] + MEM[10408];
assign MEM[19185] = MEM[4422] + MEM[7084];
assign MEM[19186] = MEM[4423] + MEM[12218];
assign MEM[19187] = MEM[4426] + MEM[5718];
assign MEM[19188] = MEM[4428] + MEM[6555];
assign MEM[19189] = MEM[4430] + MEM[6354];
assign MEM[19190] = MEM[4431] + MEM[5315];
assign MEM[19191] = MEM[4435] + MEM[4877];
assign MEM[19192] = MEM[4436] + MEM[5219];
assign MEM[19193] = MEM[4437] + MEM[6237];
assign MEM[19194] = MEM[4450] + MEM[6046];
assign MEM[19195] = MEM[4452] + MEM[13175];
assign MEM[19196] = MEM[4453] + MEM[11597];
assign MEM[19197] = MEM[4454] + MEM[4773];
assign MEM[19198] = MEM[4455] + MEM[14301];
assign MEM[19199] = MEM[4459] + MEM[9519];
assign MEM[19200] = MEM[4460] + MEM[8858];
assign MEM[19201] = MEM[4462] + MEM[12710];
assign MEM[19202] = MEM[4463] + MEM[8569];
assign MEM[19203] = MEM[4467] + MEM[9790];
assign MEM[19204] = MEM[4470] + MEM[12977];
assign MEM[19205] = MEM[4478] + MEM[8278];
assign MEM[19206] = MEM[4490] + MEM[13574];
assign MEM[19207] = MEM[4492] + MEM[9254];
assign MEM[19208] = MEM[4493] + MEM[6525];
assign MEM[19209] = MEM[4495] + MEM[13376];
assign MEM[19210] = MEM[4499] + MEM[10039];
assign MEM[19211] = MEM[4502] + MEM[7968];
assign MEM[19212] = MEM[4503] + MEM[10609];
assign MEM[19213] = MEM[4506] + MEM[7468];
assign MEM[19214] = MEM[4507] + MEM[7881];
assign MEM[19215] = MEM[4518] + MEM[9022];
assign MEM[19216] = MEM[4519] + MEM[5308];
assign MEM[19217] = MEM[4523] + MEM[5967];
assign MEM[19218] = MEM[4524] + MEM[11044];
assign MEM[19219] = MEM[4526] + MEM[5479];
assign MEM[19220] = MEM[4527] + MEM[11761];
assign MEM[19221] = MEM[4532] + MEM[11978];
assign MEM[19222] = MEM[4535] + MEM[11132];
assign MEM[19223] = MEM[4539] + MEM[9100];
assign MEM[19224] = MEM[4540] + MEM[9629];
assign MEM[19225] = MEM[4543] + MEM[10073];
assign MEM[19226] = MEM[4547] + MEM[16471];
assign MEM[19227] = MEM[4555] + MEM[12440];
assign MEM[19228] = MEM[4556] + MEM[9695];
assign MEM[19229] = MEM[4559] + MEM[7854];
assign MEM[19230] = MEM[4563] + MEM[9063];
assign MEM[19231] = MEM[4564] + MEM[5677];
assign MEM[19232] = MEM[4567] + MEM[4867];
assign MEM[19233] = MEM[4570] + MEM[11938];
assign MEM[19234] = MEM[4578] + MEM[14197];
assign MEM[19235] = MEM[4581] + MEM[4935];
assign MEM[19236] = MEM[4583] + MEM[11245];
assign MEM[19237] = MEM[4587] + MEM[8487];
assign MEM[19238] = MEM[4588] + MEM[12405];
assign MEM[19239] = MEM[4589] + MEM[14413];
assign MEM[19240] = MEM[4590] + MEM[11124];
assign MEM[19241] = MEM[4594] + MEM[8340];
assign MEM[19242] = MEM[4598] + MEM[7103];
assign MEM[19243] = MEM[4603] + MEM[10325];
assign MEM[19244] = MEM[4606] + MEM[8298];
assign MEM[19245] = MEM[4607] + MEM[14980];
assign MEM[19246] = MEM[4611] + MEM[14941];
assign MEM[19247] = MEM[4612] + MEM[10140];
assign MEM[19248] = MEM[4619] + MEM[15167];
assign MEM[19249] = MEM[4622] + MEM[5526];
assign MEM[19250] = MEM[4623] + MEM[6560];
assign MEM[19251] = MEM[4628] + MEM[7294];
assign MEM[19252] = MEM[4629] + MEM[8847];
assign MEM[19253] = MEM[4630] + MEM[10081];
assign MEM[19254] = MEM[4631] + MEM[10935];
assign MEM[19255] = MEM[4637] + MEM[12376];
assign MEM[19256] = MEM[4639] + MEM[8759];
assign MEM[19257] = MEM[4643] + MEM[7572];
assign MEM[19258] = MEM[4647] + MEM[13342];
assign MEM[19259] = MEM[4652] + MEM[7393];
assign MEM[19260] = MEM[4654] + MEM[5962];
assign MEM[19261] = MEM[4660] + MEM[8125];
assign MEM[19262] = MEM[4663] + MEM[14125];
assign MEM[19263] = MEM[4667] + MEM[7435];
assign MEM[19264] = MEM[4669] + MEM[9108];
assign MEM[19265] = MEM[4671] + MEM[11686];
assign MEM[19266] = MEM[4674] + MEM[11294];
assign MEM[19267] = MEM[4675] + MEM[8425];
assign MEM[19268] = MEM[4679] + MEM[9889];
assign MEM[19269] = MEM[4687] + MEM[11642];
assign MEM[19270] = MEM[4694] + MEM[13241];
assign MEM[19271] = MEM[4702] + MEM[5357];
assign MEM[19272] = MEM[4703] + MEM[10534];
assign MEM[19273] = MEM[4709] + MEM[10342];
assign MEM[19274] = MEM[4711] + MEM[14155];
assign MEM[19275] = MEM[4719] + MEM[11304];
assign MEM[19276] = MEM[4723] + MEM[12284];
assign MEM[19277] = MEM[4724] + MEM[8258];
assign MEM[19278] = MEM[4727] + MEM[11676];
assign MEM[19279] = MEM[4734] + MEM[4782];
assign MEM[19280] = MEM[4741] + MEM[6644];
assign MEM[19281] = MEM[4742] + MEM[7031];
assign MEM[19282] = MEM[4747] + MEM[12295];
assign MEM[19283] = MEM[4748] + MEM[10850];
assign MEM[19284] = MEM[4749] + MEM[11396];
assign MEM[19285] = MEM[4751] + MEM[10694];
assign MEM[19286] = MEM[4754] + MEM[5983];
assign MEM[19287] = MEM[4755] + MEM[12116];
assign MEM[19288] = MEM[4756] + MEM[7109];
assign MEM[19289] = MEM[4759] + MEM[12460];
assign MEM[19290] = MEM[4762] + MEM[12638];
assign MEM[19291] = MEM[4764] + MEM[8364];
assign MEM[19292] = MEM[4774] + MEM[8327];
assign MEM[19293] = MEM[4775] + MEM[4803];
assign MEM[19294] = MEM[4778] + MEM[12979];
assign MEM[19295] = MEM[4781] + MEM[9174];
assign MEM[19296] = MEM[4783] + MEM[6546];
assign MEM[19297] = MEM[4788] + MEM[12851];
assign MEM[19298] = MEM[4789] + MEM[5076];
assign MEM[19299] = MEM[4790] + MEM[5869];
assign MEM[19300] = MEM[4791] + MEM[10617];
assign MEM[19301] = MEM[4795] + MEM[11545];
assign MEM[19302] = MEM[4797] + MEM[6108];
assign MEM[19303] = MEM[4798] + MEM[7620];
assign MEM[19304] = MEM[4802] + MEM[12815];
assign MEM[19305] = MEM[4804] + MEM[5398];
assign MEM[19306] = MEM[4806] + MEM[9665];
assign MEM[19307] = MEM[4807] + MEM[5868];
assign MEM[19308] = MEM[4810] + MEM[5187];
assign MEM[19309] = MEM[4811] + MEM[9853];
assign MEM[19310] = MEM[4815] + MEM[9402];
assign MEM[19311] = MEM[4818] + MEM[12154];
assign MEM[19312] = MEM[4820] + MEM[8447];
assign MEM[19313] = MEM[4823] + MEM[12334];
assign MEM[19314] = MEM[4827] + MEM[8192];
assign MEM[19315] = MEM[4828] + MEM[5439];
assign MEM[19316] = MEM[4830] + MEM[6443];
assign MEM[19317] = MEM[4837] + MEM[7691];
assign MEM[19318] = MEM[4842] + MEM[8238];
assign MEM[19319] = MEM[4844] + MEM[8232];
assign MEM[19320] = MEM[4845] + MEM[4958];
assign MEM[19321] = MEM[4847] + MEM[5478];
assign MEM[19322] = MEM[4852] + MEM[5955];
assign MEM[19323] = MEM[4853] + MEM[9838];
assign MEM[19324] = MEM[4855] + MEM[10922];
assign MEM[19325] = MEM[4860] + MEM[12485];
assign MEM[19326] = MEM[4861] + MEM[5206];
assign MEM[19327] = MEM[4863] + MEM[14101];
assign MEM[19328] = MEM[4878] + MEM[8617];
assign MEM[19329] = MEM[4879] + MEM[10297];
assign MEM[19330] = MEM[4882] + MEM[12612];
assign MEM[19331] = MEM[4884] + MEM[6987];
assign MEM[19332] = MEM[4885] + MEM[13216];
assign MEM[19333] = MEM[4890] + MEM[10238];
assign MEM[19334] = MEM[4891] + MEM[6903];
assign MEM[19335] = MEM[4893] + MEM[12350];
assign MEM[19336] = MEM[4898] + MEM[8650];
assign MEM[19337] = MEM[4899] + MEM[8820];
assign MEM[19338] = MEM[4900] + MEM[9575];
assign MEM[19339] = MEM[4901] + MEM[5999];
assign MEM[19340] = MEM[4907] + MEM[13309];
assign MEM[19341] = MEM[4908] + MEM[13128];
assign MEM[19342] = MEM[4919] + MEM[12498];
assign MEM[19343] = MEM[4933] + MEM[9808];
assign MEM[19344] = MEM[4934] + MEM[7003];
assign MEM[19345] = MEM[4941] + MEM[13882];
assign MEM[19346] = MEM[4942] + MEM[13911];
assign MEM[19347] = MEM[4943] + MEM[12611];
assign MEM[19348] = MEM[4954] + MEM[14854];
assign MEM[19349] = MEM[4955] + MEM[13024];
assign MEM[19350] = MEM[4957] + MEM[17021];
assign MEM[19351] = MEM[4959] + MEM[13439];
assign MEM[19352] = MEM[4963] + MEM[17425];
assign MEM[19353] = MEM[4966] + MEM[6481];
assign MEM[19354] = MEM[4970] + MEM[7096];
assign MEM[19355] = MEM[4975] + MEM[8467];
assign MEM[19356] = MEM[4978] + MEM[7908];
assign MEM[19357] = MEM[4980] + MEM[15320];
assign MEM[19358] = MEM[4981] + MEM[8070];
assign MEM[19359] = MEM[4983] + MEM[8018];
assign MEM[19360] = MEM[4988] + MEM[8324];
assign MEM[19361] = MEM[4990] + MEM[10393];
assign MEM[19362] = MEM[4991] + MEM[8681];
assign MEM[19363] = MEM[4994] + MEM[8615];
assign MEM[19364] = MEM[4995] + MEM[14285];
assign MEM[19365] = MEM[5004] + MEM[13725];
assign MEM[19366] = MEM[5006] + MEM[7949];
assign MEM[19367] = MEM[5011] + MEM[12813];
assign MEM[19368] = MEM[5012] + MEM[12766];
assign MEM[19369] = MEM[5014] + MEM[13008];
assign MEM[19370] = MEM[5020] + MEM[6418];
assign MEM[19371] = MEM[5022] + MEM[8795];
assign MEM[19372] = MEM[5028] + MEM[8221];
assign MEM[19373] = MEM[5030] + MEM[15033];
assign MEM[19374] = MEM[5035] + MEM[12772];
assign MEM[19375] = MEM[5036] + MEM[10495];
assign MEM[19376] = MEM[5038] + MEM[5838];
assign MEM[19377] = MEM[5042] + MEM[13086];
assign MEM[19378] = MEM[5045] + MEM[9290];
assign MEM[19379] = MEM[5046] + MEM[7868];
assign MEM[19380] = MEM[5047] + MEM[5266];
assign MEM[19381] = MEM[5052] + MEM[16469];
assign MEM[19382] = MEM[5054] + MEM[8455];
assign MEM[19383] = MEM[5059] + MEM[7674];
assign MEM[19384] = MEM[5061] + MEM[13656];
assign MEM[19385] = MEM[5063] + MEM[8165];
assign MEM[19386] = MEM[5078] + MEM[12686];
assign MEM[19387] = MEM[5079] + MEM[10187];
assign MEM[19388] = MEM[5082] + MEM[8024];
assign MEM[19389] = MEM[5085] + MEM[9745];
assign MEM[19390] = MEM[5086] + MEM[14056];
assign MEM[19391] = MEM[5093] + MEM[11722];
assign MEM[19392] = MEM[5095] + MEM[13115];
assign MEM[19393] = MEM[5099] + MEM[12185];
assign MEM[19394] = MEM[5100] + MEM[12242];
assign MEM[19395] = MEM[5103] + MEM[8933];
assign MEM[19396] = MEM[5106] + MEM[7873];
assign MEM[19397] = MEM[5108] + MEM[13193];
assign MEM[19398] = MEM[5109] + MEM[8486];
assign MEM[19399] = MEM[5123] + MEM[8261];
assign MEM[19400] = MEM[5124] + MEM[7060];
assign MEM[19401] = MEM[5126] + MEM[11469];
assign MEM[19402] = MEM[5127] + MEM[5227];
assign MEM[19403] = MEM[5131] + MEM[14564];
assign MEM[19404] = MEM[5132] + MEM[5167];
assign MEM[19405] = MEM[5139] + MEM[12157];
assign MEM[19406] = MEM[5143] + MEM[8548];
assign MEM[19407] = MEM[5149] + MEM[6284];
assign MEM[19408] = MEM[5151] + MEM[11228];
assign MEM[19409] = MEM[5157] + MEM[7772];
assign MEM[19410] = MEM[5171] + MEM[8391];
assign MEM[19411] = MEM[5174] + MEM[7783];
assign MEM[19412] = MEM[5180] + MEM[9920];
assign MEM[19413] = MEM[5181] + MEM[7345];
assign MEM[19414] = MEM[5183] + MEM[5663];
assign MEM[19415] = MEM[5186] + MEM[12029];
assign MEM[19416] = MEM[5188] + MEM[6943];
assign MEM[19417] = MEM[5197] + MEM[8429];
assign MEM[19418] = MEM[5204] + MEM[14703];
assign MEM[19419] = MEM[5210] + MEM[12799];
assign MEM[19420] = MEM[5211] + MEM[12220];
assign MEM[19421] = MEM[5214] + MEM[7608];
assign MEM[19422] = MEM[5218] + MEM[13300];
assign MEM[19423] = MEM[5220] + MEM[12748];
assign MEM[19424] = MEM[5221] + MEM[19021];
assign MEM[19425] = MEM[5223] + MEM[10299];
assign MEM[19426] = MEM[5226] + MEM[15227];
assign MEM[19427] = MEM[5229] + MEM[9634];
assign MEM[19428] = MEM[5235] + MEM[9175];
assign MEM[19429] = MEM[5236] + MEM[10986];
assign MEM[19430] = MEM[5237] + MEM[12404];
assign MEM[19431] = MEM[5243] + MEM[5251];
assign MEM[19432] = MEM[5246] + MEM[15979];
assign MEM[19433] = MEM[5247] + MEM[5412];
assign MEM[19434] = MEM[5252] + MEM[5614];
assign MEM[19435] = MEM[5254] + MEM[10946];
assign MEM[19436] = MEM[5255] + MEM[9847];
assign MEM[19437] = MEM[5260] + MEM[5515];
assign MEM[19438] = MEM[5261] + MEM[6648];
assign MEM[19439] = MEM[5267] + MEM[9702];
assign MEM[19440] = MEM[5269] + MEM[5283];
assign MEM[19441] = MEM[5270] + MEM[6439];
assign MEM[19442] = MEM[5275] + MEM[16162];
assign MEM[19443] = MEM[5278] + MEM[9625];
assign MEM[19444] = MEM[5279] + MEM[8514];
assign MEM[19445] = MEM[5282] + MEM[13044];
assign MEM[19446] = MEM[5284] + MEM[10689];
assign MEM[19447] = MEM[5286] + MEM[6691];
assign MEM[19448] = MEM[5287] + MEM[8806];
assign MEM[19449] = MEM[5290] + MEM[7343];
assign MEM[19450] = MEM[5291] + MEM[8264];
assign MEM[19451] = MEM[5292] + MEM[10577];
assign MEM[19452] = MEM[5293] + MEM[8143];
assign MEM[19453] = MEM[5294] + MEM[8071];
assign MEM[19454] = MEM[5300] + MEM[13487];
assign MEM[19455] = MEM[5303] + MEM[9008];
assign MEM[19456] = MEM[5306] + MEM[6593];
assign MEM[19457] = MEM[5307] + MEM[11021];
assign MEM[19458] = MEM[5310] + MEM[7750];
assign MEM[19459] = MEM[5314] + MEM[6700];
assign MEM[19460] = MEM[5317] + MEM[8909];
assign MEM[19461] = MEM[5318] + MEM[12087];
assign MEM[19462] = MEM[5322] + MEM[9499];
assign MEM[19463] = MEM[5324] + MEM[7843];
assign MEM[19464] = MEM[5327] + MEM[6279];
assign MEM[19465] = MEM[5330] + MEM[10379];
assign MEM[19466] = MEM[5331] + MEM[6519];
assign MEM[19467] = MEM[5342] + MEM[11247];
assign MEM[19468] = MEM[5347] + MEM[7984];
assign MEM[19469] = MEM[5348] + MEM[8545];
assign MEM[19470] = MEM[5349] + MEM[14468];
assign MEM[19471] = MEM[5350] + MEM[11075];
assign MEM[19472] = MEM[5351] + MEM[9667];
assign MEM[19473] = MEM[5355] + MEM[11052];
assign MEM[19474] = MEM[5382] + MEM[7661];
assign MEM[19475] = MEM[5383] + MEM[12983];
assign MEM[19476] = MEM[5395] + MEM[8362];
assign MEM[19477] = MEM[5399] + MEM[6907];
assign MEM[19478] = MEM[5403] + MEM[8935];
assign MEM[19479] = MEM[5404] + MEM[6358];
assign MEM[19480] = MEM[5405] + MEM[6841];
assign MEM[19481] = MEM[5407] + MEM[11498];
assign MEM[19482] = MEM[5410] + MEM[15034];
assign MEM[19483] = MEM[5411] + MEM[5727];
assign MEM[19484] = MEM[5414] + MEM[8871];
assign MEM[19485] = MEM[5418] + MEM[6968];
assign MEM[19486] = MEM[5421] + MEM[13167];
assign MEM[19487] = MEM[5427] + MEM[6338];
assign MEM[19488] = MEM[5428] + MEM[15507];
assign MEM[19489] = MEM[5430] + MEM[11027];
assign MEM[19490] = MEM[5434] + MEM[6069];
assign MEM[19491] = MEM[5435] + MEM[10701];
assign MEM[19492] = MEM[5436] + MEM[8595];
assign MEM[19493] = MEM[5438] + MEM[6505];
assign MEM[19494] = MEM[5442] + MEM[9903];
assign MEM[19495] = MEM[5445] + MEM[12341];
assign MEM[19496] = MEM[5450] + MEM[5874];
assign MEM[19497] = MEM[5451] + MEM[9312];
assign MEM[19498] = MEM[5460] + MEM[8136];
assign MEM[19499] = MEM[5462] + MEM[13240];
assign MEM[19500] = MEM[5463] + MEM[8669];
assign MEM[19501] = MEM[5467] + MEM[12936];
assign MEM[19502] = MEM[5471] + MEM[5748];
assign MEM[19503] = MEM[5483] + MEM[8145];
assign MEM[19504] = MEM[5486] + MEM[10534];
assign MEM[19505] = MEM[5492] + MEM[7429];
assign MEM[19506] = MEM[5493] + MEM[12351];
assign MEM[19507] = MEM[5498] + MEM[16810];
assign MEM[19508] = MEM[5501] + MEM[9975];
assign MEM[19509] = MEM[5506] + MEM[7413];
assign MEM[19510] = MEM[5507] + MEM[13164];
assign MEM[19511] = MEM[5508] + MEM[6698];
assign MEM[19512] = MEM[5514] + MEM[14638];
assign MEM[19513] = MEM[5515] + MEM[13714];
assign MEM[19514] = MEM[5516] + MEM[6870];
assign MEM[19515] = MEM[5522] + MEM[12727];
assign MEM[19516] = MEM[5525] + MEM[6423];
assign MEM[19517] = MEM[5527] + MEM[13153];
assign MEM[19518] = MEM[5532] + MEM[13322];
assign MEM[19519] = MEM[5533] + MEM[11519];
assign MEM[19520] = MEM[5534] + MEM[16206];
assign MEM[19521] = MEM[5539] + MEM[12119];
assign MEM[19522] = MEM[5540] + MEM[5862];
assign MEM[19523] = MEM[5549] + MEM[7119];
assign MEM[19524] = MEM[5551] + MEM[6611];
assign MEM[19525] = MEM[5555] + MEM[5709];
assign MEM[19526] = MEM[5557] + MEM[7246];
assign MEM[19527] = MEM[5558] + MEM[11923];
assign MEM[19528] = MEM[5559] + MEM[10559];
assign MEM[19529] = MEM[5563] + MEM[7260];
assign MEM[19530] = MEM[5570] + MEM[6633];
assign MEM[19531] = MEM[5572] + MEM[6676];
assign MEM[19532] = MEM[5573] + MEM[12929];
assign MEM[19533] = MEM[5575] + MEM[12225];
assign MEM[19534] = MEM[5580] + MEM[6273];
assign MEM[19535] = MEM[5582] + MEM[5732];
assign MEM[19536] = MEM[5583] + MEM[12592];
assign MEM[19537] = MEM[5589] + MEM[8065];
assign MEM[19538] = MEM[5590] + MEM[8709];
assign MEM[19539] = MEM[5598] + MEM[11768];
assign MEM[19540] = MEM[5605] + MEM[12768];
assign MEM[19541] = MEM[5622] + MEM[13000];
assign MEM[19542] = MEM[5623] + MEM[6295];
assign MEM[19543] = MEM[5627] + MEM[12567];
assign MEM[19544] = MEM[5628] + MEM[6485];
assign MEM[19545] = MEM[5630] + MEM[7234];
assign MEM[19546] = MEM[5636] + MEM[8022];
assign MEM[19547] = MEM[5639] + MEM[11180];
assign MEM[19548] = MEM[5642] + MEM[9805];
assign MEM[19549] = MEM[5643] + MEM[12089];
assign MEM[19550] = MEM[5646] + MEM[10915];
assign MEM[19551] = MEM[5647] + MEM[13009];
assign MEM[19552] = MEM[5651] + MEM[7420];
assign MEM[19553] = MEM[5652] + MEM[6438];
assign MEM[19554] = MEM[5654] + MEM[7597];
assign MEM[19555] = MEM[5655] + MEM[12649];
assign MEM[19556] = MEM[5659] + MEM[9656];
assign MEM[19557] = MEM[5666] + MEM[9610];
assign MEM[19558] = MEM[5675] + MEM[7711];
assign MEM[19559] = MEM[5683] + MEM[7352];
assign MEM[19560] = MEM[5686] + MEM[9488];
assign MEM[19561] = MEM[5693] + MEM[14698];
assign MEM[19562] = MEM[5694] + MEM[7105];
assign MEM[19563] = MEM[5695] + MEM[8229];
assign MEM[19564] = MEM[5700] + MEM[9929];
assign MEM[19565] = MEM[5706] + MEM[11359];
assign MEM[19566] = MEM[5715] + MEM[8433];
assign MEM[19567] = MEM[5722] + MEM[6238];
assign MEM[19568] = MEM[5723] + MEM[10435];
assign MEM[19569] = MEM[5724] + MEM[12137];
assign MEM[19570] = MEM[5725] + MEM[12476];
assign MEM[19571] = MEM[5726] + MEM[12356];
assign MEM[19572] = MEM[5730] + MEM[14936];
assign MEM[19573] = MEM[5733] + MEM[6566];
assign MEM[19574] = MEM[5737] + MEM[13847];
assign MEM[19575] = MEM[5740] + MEM[13379];
assign MEM[19576] = MEM[5741] + MEM[12657];
assign MEM[19577] = MEM[5742] + MEM[10388];
assign MEM[19578] = MEM[5743] + MEM[12987];
assign MEM[19579] = MEM[5749] + MEM[11786];
assign MEM[19580] = MEM[5751] + MEM[10789];
assign MEM[19581] = MEM[5755] + MEM[6204];
assign MEM[19582] = MEM[5762] + MEM[8377];
assign MEM[19583] = MEM[5763] + MEM[7248];
assign MEM[19584] = MEM[5773] + MEM[8103];
assign MEM[19585] = MEM[5774] + MEM[9192];
assign MEM[19586] = MEM[5779] + MEM[6950];
assign MEM[19587] = MEM[5781] + MEM[13638];
assign MEM[19588] = MEM[5783] + MEM[11178];
assign MEM[19589] = MEM[5789] + MEM[7747];
assign MEM[19590] = MEM[5790] + MEM[7749];
assign MEM[19591] = MEM[5791] + MEM[10910];
assign MEM[19592] = MEM[5797] + MEM[6951];
assign MEM[19593] = MEM[5798] + MEM[9685];
assign MEM[19594] = MEM[5805] + MEM[12645];
assign MEM[19595] = MEM[5806] + MEM[15834];
assign MEM[19596] = MEM[5822] + MEM[11321];
assign MEM[19597] = MEM[5823] + MEM[16568];
assign MEM[19598] = MEM[5830] + MEM[7928];
assign MEM[19599] = MEM[5837] + MEM[14216];
assign MEM[19600] = MEM[5855] + MEM[12375];
assign MEM[19601] = MEM[5858] + MEM[9810];
assign MEM[19602] = MEM[5863] + MEM[13178];
assign MEM[19603] = MEM[5866] + MEM[13547];
assign MEM[19604] = MEM[5867] + MEM[10529];
assign MEM[19605] = MEM[5875] + MEM[8599];
assign MEM[19606] = MEM[5876] + MEM[9049];
assign MEM[19607] = MEM[5879] + MEM[11954];
assign MEM[19608] = MEM[5882] + MEM[6695];
assign MEM[19609] = MEM[5884] + MEM[10729];
assign MEM[19610] = MEM[5885] + MEM[13160];
assign MEM[19611] = MEM[5891] + MEM[13986];
assign MEM[19612] = MEM[5892] + MEM[12296];
assign MEM[19613] = MEM[5894] + MEM[15108];
assign MEM[19614] = MEM[5895] + MEM[15795];
assign MEM[19615] = MEM[5896] + MEM[8877];
assign MEM[19616] = MEM[5897] + MEM[12670];
assign MEM[19617] = MEM[5900] + MEM[8733];
assign MEM[19618] = MEM[5902] + MEM[13161];
assign MEM[19619] = MEM[5905] + MEM[9628];
assign MEM[19620] = MEM[5906] + MEM[10204];
assign MEM[19621] = MEM[5908] + MEM[13904];
assign MEM[19622] = MEM[5909] + MEM[16584];
assign MEM[19623] = MEM[5914] + MEM[8535];
assign MEM[19624] = MEM[5922] + MEM[15745];
assign MEM[19625] = MEM[5924] + MEM[11771];
assign MEM[19626] = MEM[5925] + MEM[15900];
assign MEM[19627] = MEM[5928] + MEM[14702];
assign MEM[19628] = MEM[5929] + MEM[9288];
assign MEM[19629] = MEM[5930] + MEM[7102];
assign MEM[19630] = MEM[5931] + MEM[11689];
assign MEM[19631] = MEM[5932] + MEM[12662];
assign MEM[19632] = MEM[5933] + MEM[14175];
assign MEM[19633] = MEM[5935] + MEM[14685];
assign MEM[19634] = MEM[5939] + MEM[13060];
assign MEM[19635] = MEM[5949] + MEM[7495];
assign MEM[19636] = MEM[5954] + MEM[9160];
assign MEM[19637] = MEM[5956] + MEM[8850];
assign MEM[19638] = MEM[5959] + MEM[8016];
assign MEM[19639] = MEM[5963] + MEM[8571];
assign MEM[19640] = MEM[5964] + MEM[9052];
assign MEM[19641] = MEM[5965] + MEM[10209];
assign MEM[19642] = MEM[5972] + MEM[6798];
assign MEM[19643] = MEM[5975] + MEM[12938];
assign MEM[19644] = MEM[5980] + MEM[9068];
assign MEM[19645] = MEM[5982] + MEM[7287];
assign MEM[19646] = MEM[5987] + MEM[12971];
assign MEM[19647] = MEM[5994] + MEM[8682];
assign MEM[19648] = MEM[5995] + MEM[7730];
assign MEM[19649] = MEM[6002] + MEM[13400];
assign MEM[19650] = MEM[6004] + MEM[8793];
assign MEM[19651] = MEM[6013] + MEM[7065];
assign MEM[19652] = MEM[6021] + MEM[8254];
assign MEM[19653] = MEM[6030] + MEM[7094];
assign MEM[19654] = MEM[6038] + MEM[8072];
assign MEM[19655] = MEM[6039] + MEM[3079];
assign MEM[19656] = MEM[6045] + MEM[8713];
assign MEM[19657] = MEM[6053] + MEM[13165];
assign MEM[19658] = MEM[6063] + MEM[9219];
assign MEM[19659] = MEM[6070] + MEM[8716];
assign MEM[19660] = MEM[6071] + MEM[11356];
assign MEM[19661] = MEM[6079] + MEM[13653];
assign MEM[19662] = MEM[6085] + MEM[15321];
assign MEM[19663] = MEM[6087] + MEM[6995];
assign MEM[19664] = MEM[6093] + MEM[10292];
assign MEM[19665] = MEM[6103] + MEM[11547];
assign MEM[19666] = MEM[6116] + MEM[8955];
assign MEM[19667] = MEM[6126] + MEM[7110];
assign MEM[19668] = MEM[6134] + MEM[12599];
assign MEM[19669] = MEM[6140] + MEM[13428];
assign MEM[19670] = MEM[6148] + MEM[16086];
assign MEM[19671] = MEM[6149] + MEM[7671];
assign MEM[19672] = MEM[6151] + MEM[7609];
assign MEM[19673] = MEM[6154] + MEM[12758];
assign MEM[19674] = MEM[6156] + MEM[7568];
assign MEM[19675] = MEM[6157] + MEM[8552];
assign MEM[19676] = MEM[6158] + MEM[6674];
assign MEM[19677] = MEM[6159] + MEM[12016];
assign MEM[19678] = MEM[6163] + MEM[6348];
assign MEM[19679] = MEM[6173] + MEM[11158];
assign MEM[19680] = MEM[6174] + MEM[7508];
assign MEM[19681] = MEM[6178] + MEM[8613];
assign MEM[19682] = MEM[6180] + MEM[13886];
assign MEM[19683] = MEM[6183] + MEM[12525];
assign MEM[19684] = MEM[6187] + MEM[8611];
assign MEM[19685] = MEM[6190] + MEM[7384];
assign MEM[19686] = MEM[6191] + MEM[7395];
assign MEM[19687] = MEM[6195] + MEM[8381];
assign MEM[19688] = MEM[6199] + MEM[8200];
assign MEM[19689] = MEM[6205] + MEM[7982];
assign MEM[19690] = MEM[6205] + MEM[15165];
assign MEM[19691] = MEM[6207] + MEM[15424];
assign MEM[19692] = MEM[6214] + MEM[8041];
assign MEM[19693] = MEM[6221] + MEM[8741];
assign MEM[19694] = MEM[6229] + MEM[8476];
assign MEM[19695] = MEM[6230] + MEM[8442];
assign MEM[19696] = MEM[6231] + MEM[9080];
assign MEM[19697] = MEM[6253] + MEM[7236];
assign MEM[19698] = MEM[6261] + MEM[8262];
assign MEM[19699] = MEM[6275] + MEM[9594];
assign MEM[19700] = MEM[6277] + MEM[11846];
assign MEM[19701] = MEM[6281] + MEM[12278];
assign MEM[19702] = MEM[6282] + MEM[7718];
assign MEM[19703] = MEM[6283] + MEM[7365];
assign MEM[19704] = MEM[6285] + MEM[16631];
assign MEM[19705] = MEM[6286] + MEM[11579];
assign MEM[19706] = MEM[6289] + MEM[14416];
assign MEM[19707] = MEM[6293] + MEM[6331];
assign MEM[19708] = MEM[6299] + MEM[16069];
assign MEM[19709] = MEM[6301] + MEM[13221];
assign MEM[19710] = MEM[6303] + MEM[12080];
assign MEM[19711] = MEM[6304] + MEM[15630];
assign MEM[19712] = MEM[6306] + MEM[8001];
assign MEM[19713] = MEM[6310] + MEM[13604];
assign MEM[19714] = MEM[6311] + MEM[11089];
assign MEM[19715] = MEM[6314] + MEM[16384];
assign MEM[19716] = MEM[6315] + MEM[13733];
assign MEM[19717] = MEM[6317] + MEM[10904];
assign MEM[19718] = MEM[6323] + MEM[7204];
assign MEM[19719] = MEM[6325] + MEM[9047];
assign MEM[19720] = MEM[6326] + MEM[16666];
assign MEM[19721] = MEM[6327] + MEM[7824];
assign MEM[19722] = MEM[6328] + MEM[10788];
assign MEM[19723] = MEM[6332] + MEM[13808];
assign MEM[19724] = MEM[6333] + MEM[10291];
assign MEM[19725] = MEM[6335] + MEM[10127];
assign MEM[19726] = MEM[6339] + MEM[12265];
assign MEM[19727] = MEM[6340] + MEM[12238];
assign MEM[19728] = MEM[6344] + MEM[13356];
assign MEM[19729] = MEM[6345] + MEM[8409];
assign MEM[19730] = MEM[6346] + MEM[12501];
assign MEM[19731] = MEM[6347] + MEM[7310];
assign MEM[19732] = MEM[6360] + MEM[6658];
assign MEM[19733] = MEM[6362] + MEM[9278];
assign MEM[19734] = MEM[6364] + MEM[10290];
assign MEM[19735] = MEM[6366] + MEM[9093];
assign MEM[19736] = MEM[6368] + MEM[15772];
assign MEM[19737] = MEM[6369] + MEM[11779];
assign MEM[19738] = MEM[6370] + MEM[7486];
assign MEM[19739] = MEM[6371] + MEM[6832];
assign MEM[19740] = MEM[6373] + MEM[11860];
assign MEM[19741] = MEM[6375] + MEM[9409];
assign MEM[19742] = MEM[6379] + MEM[8037];
assign MEM[19743] = MEM[6381] + MEM[11577];
assign MEM[19744] = MEM[6385] + MEM[12374];
assign MEM[19745] = MEM[6389] + MEM[7686];
assign MEM[19746] = MEM[6412] + MEM[9484];
assign MEM[19747] = MEM[6414] + MEM[13836];
assign MEM[19748] = MEM[6415] + MEM[8170];
assign MEM[19749] = MEM[6416] + MEM[6568];
assign MEM[19750] = MEM[6424] + MEM[9521];
assign MEM[19751] = MEM[6426] + MEM[9330];
assign MEM[19752] = MEM[6427] + MEM[12188];
assign MEM[19753] = MEM[6430] + MEM[10324];
assign MEM[19754] = MEM[6434] + MEM[11140];
assign MEM[19755] = MEM[6435] + MEM[9210];
assign MEM[19756] = MEM[6436] + MEM[10629];
assign MEM[19757] = MEM[6440] + MEM[12336];
assign MEM[19758] = MEM[6441] + MEM[7780];
assign MEM[19759] = MEM[6462] + MEM[12454];
assign MEM[19760] = MEM[6468] + MEM[10832];
assign MEM[19761] = MEM[6471] + MEM[14417];
assign MEM[19762] = MEM[6472] + MEM[8598];
assign MEM[19763] = MEM[6474] + MEM[12931];
assign MEM[19764] = MEM[6476] + MEM[11113];
assign MEM[19765] = MEM[6477] + MEM[12106];
assign MEM[19766] = MEM[6480] + MEM[8466];
assign MEM[19767] = MEM[6488] + MEM[11160];
assign MEM[19768] = MEM[6490] + MEM[11704];
assign MEM[19769] = MEM[6491] + MEM[10632];
assign MEM[19770] = MEM[6493] + MEM[11149];
assign MEM[19771] = MEM[6495] + MEM[9072];
assign MEM[19772] = MEM[6496] + MEM[9596];
assign MEM[19773] = MEM[6499] + MEM[12168];
assign MEM[19774] = MEM[6500] + MEM[11050];
assign MEM[19775] = MEM[6501] + MEM[10007];
assign MEM[19776] = MEM[6506] + MEM[8162];
assign MEM[19777] = MEM[6507] + MEM[14085];
assign MEM[19778] = MEM[6513] + MEM[10282];
assign MEM[19779] = MEM[6524] + MEM[11877];
assign MEM[19780] = MEM[6536] + MEM[13046];
assign MEM[19781] = MEM[6547] + MEM[7903];
assign MEM[19782] = MEM[6548] + MEM[7736];
assign MEM[19783] = MEM[6556] + MEM[7734];
assign MEM[19784] = MEM[6561] + MEM[11252];
assign MEM[19785] = MEM[6563] + MEM[12172];
assign MEM[19786] = MEM[6565] + MEM[13084];
assign MEM[19787] = MEM[6567] + MEM[11290];
assign MEM[19788] = MEM[6576] + MEM[13136];
assign MEM[19789] = MEM[6577] + MEM[13788];
assign MEM[19790] = MEM[6581] + MEM[14750];
assign MEM[19791] = MEM[6588] + MEM[8586];
assign MEM[19792] = MEM[6589] + MEM[8925];
assign MEM[19793] = MEM[6590] + MEM[10734];
assign MEM[19794] = MEM[6605] + MEM[13860];
assign MEM[19795] = MEM[6608] + MEM[7548];
assign MEM[19796] = MEM[6609] + MEM[12865];
assign MEM[19797] = MEM[6616] + MEM[8490];
assign MEM[19798] = MEM[6616] + MEM[9606];
assign MEM[19799] = MEM[6620] + MEM[8194];
assign MEM[19800] = MEM[6631] + MEM[12086];
assign MEM[19801] = MEM[6649] + MEM[12804];
assign MEM[19802] = MEM[6656] + MEM[8892];
assign MEM[19803] = MEM[6657] + MEM[7485];
assign MEM[19804] = MEM[6659] + MEM[8916];
assign MEM[19805] = MEM[6661] + MEM[7788];
assign MEM[19806] = MEM[6663] + MEM[9614];
assign MEM[19807] = MEM[6668] + MEM[13209];
assign MEM[19808] = MEM[6672] + MEM[12510];
assign MEM[19809] = MEM[6673] + MEM[7350];
assign MEM[19810] = MEM[6675] + MEM[10634];
assign MEM[19811] = MEM[6678] + MEM[13861];
assign MEM[19812] = MEM[6681] + MEM[12402];
assign MEM[19813] = MEM[6682] + MEM[9385];
assign MEM[19814] = MEM[6685] + MEM[13757];
assign MEM[19815] = MEM[6692] + MEM[17087];
assign MEM[19816] = MEM[6693] + MEM[13756];
assign MEM[19817] = MEM[6694] + MEM[17707];
assign MEM[19818] = MEM[6696] + MEM[12408];
assign MEM[19819] = MEM[6701] + MEM[10786];
assign MEM[19820] = MEM[6702] + MEM[7731];
assign MEM[19821] = MEM[6705] + MEM[12034];
assign MEM[19822] = MEM[6716] + MEM[7269];
assign MEM[19823] = MEM[6736] + MEM[6981];
assign MEM[19824] = MEM[6738] + MEM[11925];
assign MEM[19825] = MEM[6741] + MEM[13000];
assign MEM[19826] = MEM[6742] + MEM[14061];
assign MEM[19827] = MEM[6745] + MEM[10139];
assign MEM[19828] = MEM[6748] + MEM[8248];
assign MEM[19829] = MEM[6749] + MEM[11014];
assign MEM[19830] = MEM[6750] + MEM[9380];
assign MEM[19831] = MEM[6751] + MEM[12078];
assign MEM[19832] = MEM[6752] + MEM[8167];
assign MEM[19833] = MEM[6754] + MEM[6996];
assign MEM[19834] = MEM[6774] + MEM[7910];
assign MEM[19835] = MEM[6775] + MEM[13826];
assign MEM[19836] = MEM[6785] + MEM[7209];
assign MEM[19837] = MEM[6787] + MEM[8559];
assign MEM[19838] = MEM[6795] + MEM[9165];
assign MEM[19839] = MEM[6796] + MEM[9270];
assign MEM[19840] = MEM[6799] + MEM[12360];
assign MEM[19841] = MEM[6802] + MEM[12247];
assign MEM[19842] = MEM[6805] + MEM[8782];
assign MEM[19843] = MEM[6809] + MEM[12709];
assign MEM[19844] = MEM[6814] + MEM[11139];
assign MEM[19845] = MEM[6815] + MEM[15203];
assign MEM[19846] = MEM[6816] + MEM[9382];
assign MEM[19847] = MEM[6817] + MEM[9283];
assign MEM[19848] = MEM[6819] + MEM[9166];
assign MEM[19849] = MEM[6820] + MEM[10847];
assign MEM[19850] = MEM[6827] + MEM[13237];
assign MEM[19851] = MEM[6828] + MEM[12747];
assign MEM[19852] = MEM[6831] + MEM[9328];
assign MEM[19853] = MEM[6836] + MEM[10487];
assign MEM[19854] = MEM[6844] + MEM[8689];
assign MEM[19855] = MEM[6845] + MEM[14115];
assign MEM[19856] = MEM[6848] + MEM[6921];
assign MEM[19857] = MEM[6849] + MEM[10902];
assign MEM[19858] = MEM[6859] + MEM[8747];
assign MEM[19859] = MEM[6871] + MEM[8579];
assign MEM[19860] = MEM[6872] + MEM[14279];
assign MEM[19861] = MEM[6874] + MEM[8414];
assign MEM[19862] = MEM[6877] + MEM[9342];
assign MEM[19863] = MEM[6879] + MEM[8121];
assign MEM[19864] = MEM[6880] + MEM[6938];
assign MEM[19865] = MEM[6886] + MEM[13198];
assign MEM[19866] = MEM[6889] + MEM[7664];
assign MEM[19867] = MEM[6896] + MEM[7245];
assign MEM[19868] = MEM[6899] + MEM[7562];
assign MEM[19869] = MEM[6900] + MEM[7619];
assign MEM[19870] = MEM[6910] + MEM[8649];
assign MEM[19871] = MEM[6915] + MEM[12452];
assign MEM[19872] = MEM[6916] + MEM[15020];
assign MEM[19873] = MEM[6924] + MEM[14448];
assign MEM[19874] = MEM[6931] + MEM[15110];
assign MEM[19875] = MEM[6932] + MEM[15010];
assign MEM[19876] = MEM[6939] + MEM[7569];
assign MEM[19877] = MEM[6940] + MEM[11046];
assign MEM[19878] = MEM[6944] + MEM[12463];
assign MEM[19879] = MEM[6947] + MEM[11468];
assign MEM[19880] = MEM[6948] + MEM[8810];
assign MEM[19881] = MEM[6949] + MEM[12026];
assign MEM[19882] = MEM[6952] + MEM[12819];
assign MEM[19883] = MEM[6957] + MEM[12617];
assign MEM[19884] = MEM[6958] + MEM[12791];
assign MEM[19885] = MEM[6960] + MEM[9994];
assign MEM[19886] = MEM[6965] + MEM[7459];
assign MEM[19887] = MEM[6967] + MEM[12262];
assign MEM[19888] = MEM[6970] + MEM[14454];
assign MEM[19889] = MEM[6971] + MEM[15542];
assign MEM[19890] = MEM[6977] + MEM[13442];
assign MEM[19891] = MEM[6983] + MEM[11479];
assign MEM[19892] = MEM[6984] + MEM[11403];
assign MEM[19893] = MEM[6985] + MEM[7683];
assign MEM[19894] = MEM[6994] + MEM[13687];
assign MEM[19895] = MEM[6997] + MEM[14745];
assign MEM[19896] = MEM[6998] + MEM[13837];
assign MEM[19897] = MEM[6999] + MEM[9977];
assign MEM[19898] = MEM[7000] + MEM[8046];
assign MEM[19899] = MEM[7001] + MEM[8315];
assign MEM[19900] = MEM[7011] + MEM[9746];
assign MEM[19901] = MEM[7013] + MEM[12286];
assign MEM[19902] = MEM[7016] + MEM[12385];
assign MEM[19903] = MEM[7018] + MEM[12677];
assign MEM[19904] = MEM[7019] + MEM[8811];
assign MEM[19905] = MEM[7020] + MEM[14472];
assign MEM[19906] = MEM[7022] + MEM[10878];
assign MEM[19907] = MEM[7023] + MEM[8882];
assign MEM[19908] = MEM[7026] + MEM[8385];
assign MEM[19909] = MEM[7028] + MEM[12196];
assign MEM[19910] = MEM[7033] + MEM[13893];
assign MEM[19911] = MEM[7037] + MEM[8632];
assign MEM[19912] = MEM[7039] + MEM[15128];
assign MEM[19913] = MEM[7040] + MEM[14758];
assign MEM[19914] = MEM[7041] + MEM[10795];
assign MEM[19915] = MEM[7046] + MEM[14805];
assign MEM[19916] = MEM[7051] + MEM[12729];
assign MEM[19917] = MEM[7052] + MEM[7431];
assign MEM[19918] = MEM[7053] + MEM[9708];
assign MEM[19919] = MEM[7054] + MEM[12161];
assign MEM[19920] = MEM[7056] + MEM[7419];
assign MEM[19921] = MEM[7058] + MEM[12893];
assign MEM[19922] = MEM[7061] + MEM[13007];
assign MEM[19923] = MEM[7062] + MEM[9003];
assign MEM[19924] = MEM[7063] + MEM[8849];
assign MEM[19925] = MEM[7069] + MEM[14210];
assign MEM[19926] = MEM[7076] + MEM[9460];
assign MEM[19927] = MEM[7083] + MEM[8765];
assign MEM[19928] = MEM[7085] + MEM[9646];
assign MEM[19929] = MEM[7087] + MEM[9397];
assign MEM[19930] = MEM[7089] + MEM[8344];
assign MEM[19931] = MEM[7098] + MEM[8393];
assign MEM[19932] = MEM[7099] + MEM[10941];
assign MEM[19933] = MEM[7100] + MEM[15254];
assign MEM[19934] = MEM[7101] + MEM[13868];
assign MEM[19935] = MEM[7106] + MEM[9755];
assign MEM[19936] = MEM[7107] + MEM[8678];
assign MEM[19937] = MEM[7114] + MEM[13179];
assign MEM[19938] = MEM[7116] + MEM[14669];
assign MEM[19939] = MEM[7118] + MEM[8770];
assign MEM[19940] = MEM[7121] + MEM[9573];
assign MEM[19941] = MEM[7126] + MEM[7732];
assign MEM[19942] = MEM[7129] + MEM[8602];
assign MEM[19943] = MEM[7133] + MEM[9001];
assign MEM[19944] = MEM[7134] + MEM[15072];
assign MEM[19945] = MEM[7139] + MEM[10244];
assign MEM[19946] = MEM[7140] + MEM[12254];
assign MEM[19947] = MEM[7141] + MEM[7706];
assign MEM[19948] = MEM[7144] + MEM[11379];
assign MEM[19949] = MEM[7148] + MEM[7993];
assign MEM[19950] = MEM[7154] + MEM[8943];
assign MEM[19951] = MEM[7155] + MEM[14209];
assign MEM[19952] = MEM[7159] + MEM[9979];
assign MEM[19953] = MEM[7160] + MEM[8068];
assign MEM[19954] = MEM[7161] + MEM[11714];
assign MEM[19955] = MEM[7162] + MEM[12298];
assign MEM[19956] = MEM[7169] + MEM[12842];
assign MEM[19957] = MEM[7170] + MEM[12480];
assign MEM[19958] = MEM[7171] + MEM[12920];
assign MEM[19959] = MEM[7172] + MEM[8977];
assign MEM[19960] = MEM[7173] + MEM[11746];
assign MEM[19961] = MEM[7175] + MEM[7377];
assign MEM[19962] = MEM[7176] + MEM[12271];
assign MEM[19963] = MEM[7184] + MEM[14020];
assign MEM[19964] = MEM[7197] + MEM[12771];
assign MEM[19965] = MEM[7199] + MEM[10613];
assign MEM[19966] = MEM[7200] + MEM[15043];
assign MEM[19967] = MEM[7201] + MEM[12269];
assign MEM[19968] = MEM[7202] + MEM[7378];
assign MEM[19969] = MEM[7206] + MEM[11623];
assign MEM[19970] = MEM[7213] + MEM[10163];
assign MEM[19971] = MEM[7216] + MEM[8333];
assign MEM[19972] = MEM[7219] + MEM[8619];
assign MEM[19973] = MEM[7224] + MEM[10708];
assign MEM[19974] = MEM[7237] + MEM[7930];
assign MEM[19975] = MEM[7239] + MEM[14951];
assign MEM[19976] = MEM[7241] + MEM[13746];
assign MEM[19977] = MEM[7242] + MEM[12666];
assign MEM[19978] = MEM[7244] + MEM[10002];
assign MEM[19979] = MEM[7249] + MEM[8415];
assign MEM[19980] = MEM[7252] + MEM[12398];
assign MEM[19981] = MEM[7254] + MEM[11242];
assign MEM[19982] = MEM[7257] + MEM[13256];
assign MEM[19983] = MEM[7261] + MEM[8179];
assign MEM[19984] = MEM[7268] + MEM[8239];
assign MEM[19985] = MEM[7270] + MEM[13864];
assign MEM[19986] = MEM[7272] + MEM[17476];
assign MEM[19987] = MEM[7274] + MEM[12232];
assign MEM[19988] = MEM[7276] + MEM[11203];
assign MEM[19989] = MEM[7277] + MEM[11071];
assign MEM[19990] = MEM[7278] + MEM[14267];
assign MEM[19991] = MEM[7280] + MEM[12786];
assign MEM[19992] = MEM[7288] + MEM[12331];
assign MEM[19993] = MEM[7293] + MEM[13431];
assign MEM[19994] = MEM[7298] + MEM[8015];
assign MEM[19995] = MEM[7299] + MEM[9276];
assign MEM[19996] = MEM[7300] + MEM[8276];
assign MEM[19997] = MEM[7301] + MEM[9611];
assign MEM[19998] = MEM[7302] + MEM[12478];
assign MEM[19999] = MEM[7306] + MEM[12400];
assign MEM[20000] = MEM[7311] + MEM[11684];
assign MEM[20001] = MEM[7312] + MEM[13244];
assign MEM[20002] = MEM[7316] + MEM[8621];
assign MEM[20003] = MEM[7317] + MEM[7837];
assign MEM[20004] = MEM[7321] + MEM[10722];
assign MEM[20005] = MEM[7326] + MEM[11517];
assign MEM[20006] = MEM[7327] + MEM[7454];
assign MEM[20007] = MEM[7329] + MEM[13553];
assign MEM[20008] = MEM[7335] + MEM[10686];
assign MEM[20009] = MEM[7338] + MEM[13040];
assign MEM[20010] = MEM[7339] + MEM[9234];
assign MEM[20011] = MEM[7357] + MEM[8691];
assign MEM[20012] = MEM[7358] + MEM[12447];
assign MEM[20013] = MEM[7368] + MEM[15116];
assign MEM[20014] = MEM[7371] + MEM[14015];
assign MEM[20015] = MEM[7373] + MEM[14763];
assign MEM[20016] = MEM[7375] + MEM[13749];
assign MEM[20017] = MEM[7380] + MEM[10531];
assign MEM[20018] = MEM[7381] + MEM[8737];
assign MEM[20019] = MEM[7382] + MEM[12394];
assign MEM[20020] = MEM[7387] + MEM[7838];
assign MEM[20021] = MEM[7392] + MEM[7911];
assign MEM[20022] = MEM[7403] + MEM[8332];
assign MEM[20023] = MEM[7409] + MEM[16158];
assign MEM[20024] = MEM[7411] + MEM[10779];
assign MEM[20025] = MEM[7418] + MEM[11222];
assign MEM[20026] = MEM[7422] + MEM[10633];
assign MEM[20027] = MEM[7430] + MEM[8479];
assign MEM[20028] = MEM[7432] + MEM[14309];
assign MEM[20029] = MEM[7434] + MEM[9935];
assign MEM[20030] = MEM[7439] + MEM[14712];
assign MEM[20031] = MEM[7442] + MEM[11243];
assign MEM[20032] = MEM[7445] + MEM[7842];
assign MEM[20033] = MEM[7451] + MEM[8293];
assign MEM[20034] = MEM[7457] + MEM[10944];
assign MEM[20035] = MEM[7464] + MEM[13581];
assign MEM[20036] = MEM[7470] + MEM[11720];
assign MEM[20037] = MEM[7472] + MEM[9548];
assign MEM[20038] = MEM[7480] + MEM[12627];
assign MEM[20039] = MEM[7481] + MEM[13762];
assign MEM[20040] = MEM[7482] + MEM[13952];
assign MEM[20041] = MEM[7506] + MEM[7755];
assign MEM[20042] = MEM[7507] + MEM[15482];
assign MEM[20043] = MEM[7509] + MEM[12571];
assign MEM[20044] = MEM[7511] + MEM[11407];
assign MEM[20045] = MEM[7512] + MEM[11564];
assign MEM[20046] = MEM[7518] + MEM[9867];
assign MEM[20047] = MEM[7523] + MEM[7712];
assign MEM[20048] = MEM[7529] + MEM[12869];
assign MEM[20049] = MEM[7530] + MEM[11901];
assign MEM[20050] = MEM[7536] + MEM[14211];
assign MEM[20051] = MEM[7537] + MEM[8520];
assign MEM[20052] = MEM[7538] + MEM[10893];
assign MEM[20053] = MEM[7539] + MEM[6309];
assign MEM[20054] = MEM[7545] + MEM[9540];
assign MEM[20055] = MEM[7546] + MEM[13689];
assign MEM[20056] = MEM[7552] + MEM[8130];
assign MEM[20057] = MEM[7559] + MEM[8843];
assign MEM[20058] = MEM[7567] + MEM[8271];
assign MEM[20059] = MEM[7570] + MEM[11583];
assign MEM[20060] = MEM[7571] + MEM[11048];
assign MEM[20061] = MEM[7573] + MEM[13743];
assign MEM[20062] = MEM[7590] + MEM[9619];
assign MEM[20063] = MEM[7592] + MEM[12852];
assign MEM[20064] = MEM[7593] + MEM[13092];
assign MEM[20065] = MEM[7596] + MEM[11006];
assign MEM[20066] = MEM[7598] + MEM[11189];
assign MEM[20067] = MEM[7599] + MEM[7678];
assign MEM[20068] = MEM[7601] + MEM[8758];
assign MEM[20069] = MEM[7602] + MEM[13692];
assign MEM[20070] = MEM[7605] + MEM[11153];
assign MEM[20071] = MEM[7606] + MEM[8457];
assign MEM[20072] = MEM[7610] + MEM[8685];
assign MEM[20073] = MEM[7611] + MEM[8577];
assign MEM[20074] = MEM[7612] + MEM[14095];
assign MEM[20075] = MEM[7613] + MEM[12092];
assign MEM[20076] = MEM[7614] + MEM[12565];
assign MEM[20077] = MEM[7618] + MEM[8056];
assign MEM[20078] = MEM[7623] + MEM[12191];
assign MEM[20079] = MEM[7624] + MEM[13764];
assign MEM[20080] = MEM[7625] + MEM[8927];
assign MEM[20081] = MEM[7627] + MEM[10591];
assign MEM[20082] = MEM[7628] + MEM[9543];
assign MEM[20083] = MEM[7631] + MEM[8246];
assign MEM[20084] = MEM[7643] + MEM[10894];
assign MEM[20085] = MEM[7645] + MEM[9825];
assign MEM[20086] = MEM[7646] + MEM[13171];
assign MEM[20087] = MEM[7649] + MEM[12555];
assign MEM[20088] = MEM[7650] + MEM[9423];
assign MEM[20089] = MEM[7651] + MEM[15769];
assign MEM[20090] = MEM[7652] + MEM[8213];
assign MEM[20091] = MEM[7654] + MEM[11560];
assign MEM[20092] = MEM[7655] + MEM[9691];
assign MEM[20093] = MEM[7657] + MEM[8537];
assign MEM[20094] = MEM[7668] + MEM[10284];
assign MEM[20095] = MEM[7669] + MEM[11195];
assign MEM[20096] = MEM[7672] + MEM[11276];
assign MEM[20097] = MEM[7675] + MEM[10964];
assign MEM[20098] = MEM[7676] + MEM[9188];
assign MEM[20099] = MEM[7679] + MEM[8277];
assign MEM[20100] = MEM[7681] + MEM[10074];
assign MEM[20101] = MEM[7684] + MEM[10042];
assign MEM[20102] = MEM[7688] + MEM[13677];
assign MEM[20103] = MEM[7690] + MEM[15077];
assign MEM[20104] = MEM[7692] + MEM[11768];
assign MEM[20105] = MEM[7694] + MEM[7728];
assign MEM[20106] = MEM[7696] + MEM[9949];
assign MEM[20107] = MEM[7699] + MEM[7710];
assign MEM[20108] = MEM[7700] + MEM[14452];
assign MEM[20109] = MEM[7701] + MEM[10956];
assign MEM[20110] = MEM[7703] + MEM[9269];
assign MEM[20111] = MEM[7704] + MEM[11585];
assign MEM[20112] = MEM[7705] + MEM[11167];
assign MEM[20113] = MEM[7708] + MEM[7851];
assign MEM[20114] = MEM[7714] + MEM[9802];
assign MEM[20115] = MEM[7716] + MEM[8176];
assign MEM[20116] = MEM[7717] + MEM[8231];
assign MEM[20117] = MEM[7719] + MEM[12079];
assign MEM[20118] = MEM[7722] + MEM[8268];
assign MEM[20119] = MEM[7725] + MEM[7878];
assign MEM[20120] = MEM[7726] + MEM[8110];
assign MEM[20121] = MEM[7729] + MEM[15006];
assign MEM[20122] = MEM[7735] + MEM[8210];
assign MEM[20123] = MEM[7739] + MEM[12544];
assign MEM[20124] = MEM[7745] + MEM[11076];
assign MEM[20125] = MEM[7757] + MEM[10454];
assign MEM[20126] = MEM[7760] + MEM[14918];
assign MEM[20127] = MEM[7773] + MEM[11260];
assign MEM[20128] = MEM[7775] + MEM[15476];
assign MEM[20129] = MEM[7778] + MEM[13062];
assign MEM[20130] = MEM[7782] + MEM[8637];
assign MEM[20131] = MEM[7784] + MEM[8722];
assign MEM[20132] = MEM[7785] + MEM[11814];
assign MEM[20133] = MEM[7786] + MEM[14636];
assign MEM[20134] = MEM[7787] + MEM[10269];
assign MEM[20135] = MEM[7794] + MEM[8112];
assign MEM[20136] = MEM[7805] + MEM[8026];
assign MEM[20137] = MEM[7808] + MEM[15032];
assign MEM[20138] = MEM[7810] + MEM[9185];
assign MEM[20139] = MEM[7811] + MEM[9141];
assign MEM[20140] = MEM[7812] + MEM[10766];
assign MEM[20141] = MEM[7819] + MEM[11619];
assign MEM[20142] = MEM[7825] + MEM[11272];
assign MEM[20143] = MEM[7827] + MEM[11007];
assign MEM[20144] = MEM[7828] + MEM[9556];
assign MEM[20145] = MEM[7835] + MEM[9415];
assign MEM[20146] = MEM[7836] + MEM[10995];
assign MEM[20147] = MEM[7839] + MEM[12872];
assign MEM[20148] = MEM[7840] + MEM[8692];
assign MEM[20149] = MEM[7845] + MEM[9337];
assign MEM[20150] = MEM[7846] + MEM[9961];
assign MEM[20151] = MEM[7852] + MEM[12348];
assign MEM[20152] = MEM[7857] + MEM[7902];
assign MEM[20153] = MEM[7860] + MEM[7871];
assign MEM[20154] = MEM[7862] + MEM[8748];
assign MEM[20155] = MEM[7864] + MEM[16294];
assign MEM[20156] = MEM[7872] + MEM[14858];
assign MEM[20157] = MEM[7874] + MEM[11079];
assign MEM[20158] = MEM[7876] + MEM[14424];
assign MEM[20159] = MEM[7882] + MEM[10996];
assign MEM[20160] = MEM[7883] + MEM[10625];
assign MEM[20161] = MEM[7889] + MEM[13022];
assign MEM[20162] = MEM[7890] + MEM[11855];
assign MEM[20163] = MEM[7891] + MEM[13401];
assign MEM[20164] = MEM[7897] + MEM[11053];
assign MEM[20165] = MEM[7901] + MEM[11734];
assign MEM[20166] = MEM[7912] + MEM[10580];
assign MEM[20167] = MEM[7913] + MEM[10371];
assign MEM[20168] = MEM[7914] + MEM[12862];
assign MEM[20169] = MEM[7918] + MEM[10200];
assign MEM[20170] = MEM[7919] + MEM[13646];
assign MEM[20171] = MEM[7922] + MEM[13367];
assign MEM[20172] = MEM[7924] + MEM[13003];
assign MEM[20173] = MEM[7925] + MEM[8953];
assign MEM[20174] = MEM[7926] + MEM[12590];
assign MEM[20175] = MEM[7927] + MEM[6155];
assign MEM[20176] = MEM[7932] + MEM[12504];
assign MEM[20177] = MEM[7938] + MEM[8677];
assign MEM[20178] = MEM[7942] + MEM[11590];
assign MEM[20179] = MEM[7944] + MEM[15292];
assign MEM[20180] = MEM[7948] + MEM[10180];
assign MEM[20181] = MEM[7951] + MEM[9512];
assign MEM[20182] = MEM[7960] + MEM[13357];
assign MEM[20183] = MEM[7963] + MEM[13797];
assign MEM[20184] = MEM[7966] + MEM[12910];
assign MEM[20185] = MEM[7969] + MEM[12908];
assign MEM[20186] = MEM[7971] + MEM[13285];
assign MEM[20187] = MEM[7974] + MEM[12564];
assign MEM[20188] = MEM[7978] + MEM[8846];
assign MEM[20189] = MEM[7979] + MEM[14573];
assign MEM[20190] = MEM[7980] + MEM[16642];
assign MEM[20191] = MEM[7981] + MEM[8982];
assign MEM[20192] = MEM[7986] + MEM[10084];
assign MEM[20193] = MEM[7992] + MEM[12103];
assign MEM[20194] = MEM[8003] + MEM[9242];
assign MEM[20195] = MEM[8005] + MEM[10053];
assign MEM[20196] = MEM[8011] + MEM[11600];
assign MEM[20197] = MEM[8012] + MEM[9151];
assign MEM[20198] = MEM[8021] + MEM[12583];
assign MEM[20199] = MEM[8023] + MEM[10107];
assign MEM[20200] = MEM[8031] + MEM[9230];
assign MEM[20201] = MEM[8034] + MEM[13110];
assign MEM[20202] = MEM[8035] + MEM[8456];
assign MEM[20203] = MEM[8038] + MEM[8932];
assign MEM[20204] = MEM[8040] + MEM[10728];
assign MEM[20205] = MEM[8044] + MEM[8879];
assign MEM[20206] = MEM[8050] + MEM[8139];
assign MEM[20207] = MEM[8052] + MEM[9106];
assign MEM[20208] = MEM[8053] + MEM[9313];
assign MEM[20209] = MEM[8054] + MEM[9688];
assign MEM[20210] = MEM[8057] + MEM[12722];
assign MEM[20211] = MEM[8061] + MEM[11286];
assign MEM[20212] = MEM[8062] + MEM[9989];
assign MEM[20213] = MEM[8064] + MEM[9718];
assign MEM[20214] = MEM[8069] + MEM[8450];
assign MEM[20215] = MEM[8073] + MEM[8319];
assign MEM[20216] = MEM[8076] + MEM[12283];
assign MEM[20217] = MEM[8077] + MEM[13528];
assign MEM[20218] = MEM[8079] + MEM[9544];
assign MEM[20219] = MEM[8080] + MEM[8597];
assign MEM[20220] = MEM[8087] + MEM[8812];
assign MEM[20221] = MEM[8089] + MEM[12312];
assign MEM[20222] = MEM[8096] + MEM[12475];
assign MEM[20223] = MEM[8097] + MEM[8911];
assign MEM[20224] = MEM[8098] + MEM[12730];
assign MEM[20225] = MEM[8099] + MEM[14607];
assign MEM[20226] = MEM[8100] + MEM[13410];
assign MEM[20227] = MEM[8106] + MEM[13301];
assign MEM[20228] = MEM[8107] + MEM[12594];
assign MEM[20229] = MEM[8109] + MEM[11224];
assign MEM[20230] = MEM[8111] + MEM[8382];
assign MEM[20231] = MEM[8113] + MEM[8416];
assign MEM[20232] = MEM[8115] + MEM[8565];
assign MEM[20233] = MEM[8117] + MEM[10272];
assign MEM[20234] = MEM[8119] + MEM[13795];
assign MEM[20235] = MEM[8122] + MEM[11129];
assign MEM[20236] = MEM[8123] + MEM[8744];
assign MEM[20237] = MEM[8126] + MEM[13693];
assign MEM[20238] = MEM[8127] + MEM[8426];
assign MEM[20239] = MEM[8128] + MEM[12321];
assign MEM[20240] = MEM[8129] + MEM[12756];
assign MEM[20241] = MEM[8133] + MEM[10224];
assign MEM[20242] = MEM[8135] + MEM[8854];
assign MEM[20243] = MEM[8137] + MEM[13938];
assign MEM[20244] = MEM[8140] + MEM[14498];
assign MEM[20245] = MEM[8142] + MEM[9101];
assign MEM[20246] = MEM[8144] + MEM[14782];
assign MEM[20247] = MEM[8147] + MEM[10162];
assign MEM[20248] = MEM[8148] + MEM[8760];
assign MEM[20249] = MEM[8159] + MEM[13751];
assign MEM[20250] = MEM[8160] + MEM[8991];
assign MEM[20251] = MEM[8164] + MEM[8357];
assign MEM[20252] = MEM[8166] + MEM[11563];
assign MEM[20253] = MEM[8168] + MEM[11910];
assign MEM[20254] = MEM[8172] + MEM[12594];
assign MEM[20255] = MEM[8173] + MEM[13267];
assign MEM[20256] = MEM[8174] + MEM[13935];
assign MEM[20257] = MEM[8175] + MEM[9411];
assign MEM[20258] = MEM[8180] + MEM[10186];
assign MEM[20259] = MEM[8181] + MEM[10690];
assign MEM[20260] = MEM[8189] + MEM[9883];
assign MEM[20261] = MEM[8190] + MEM[8612];
assign MEM[20262] = MEM[8195] + MEM[13116];
assign MEM[20263] = MEM[8199] + MEM[9235];
assign MEM[20264] = MEM[8202] + MEM[8307];
assign MEM[20265] = MEM[8203] + MEM[9222];
assign MEM[20266] = MEM[8206] + MEM[12357];
assign MEM[20267] = MEM[8207] + MEM[8216];
assign MEM[20268] = MEM[8208] + MEM[11830];
assign MEM[20269] = MEM[8209] + MEM[11292];
assign MEM[20270] = MEM[8214] + MEM[9704];
assign MEM[20271] = MEM[8215] + MEM[8303];
assign MEM[20272] = MEM[8218] + MEM[9323];
assign MEM[20273] = MEM[8220] + MEM[12537];
assign MEM[20274] = MEM[8222] + MEM[14291];
assign MEM[20275] = MEM[8224] + MEM[13731];
assign MEM[20276] = MEM[8225] + MEM[10395];
assign MEM[20277] = MEM[8227] + MEM[12387];
assign MEM[20278] = MEM[8236] + MEM[8684];
assign MEM[20279] = MEM[8242] + MEM[13332];
assign MEM[20280] = MEM[8247] + MEM[13076];
assign MEM[20281] = MEM[8250] + MEM[8674];
assign MEM[20282] = MEM[8251] + MEM[9508];
assign MEM[20283] = MEM[8255] + MEM[9676];
assign MEM[20284] = MEM[8256] + MEM[9895];
assign MEM[20285] = MEM[8257] + MEM[10799];
assign MEM[20286] = MEM[8259] + MEM[15379];
assign MEM[20287] = MEM[8260] + MEM[12751];
assign MEM[20288] = MEM[8270] + MEM[9971];
assign MEM[20289] = MEM[8273] + MEM[9125];
assign MEM[20290] = MEM[8275] + MEM[10041];
assign MEM[20291] = MEM[8280] + MEM[13493];
assign MEM[20292] = MEM[8281] + MEM[8789];
assign MEM[20293] = MEM[8283] + MEM[13575];
assign MEM[20294] = MEM[8285] + MEM[12106];
assign MEM[20295] = MEM[8290] + MEM[12637];
assign MEM[20296] = MEM[8291] + MEM[9542];
assign MEM[20297] = MEM[8296] + MEM[11020];
assign MEM[20298] = MEM[8297] + MEM[8572];
assign MEM[20299] = MEM[8300] + MEM[13857];
assign MEM[20300] = MEM[8305] + MEM[14385];
assign MEM[20301] = MEM[8306] + MEM[10699];
assign MEM[20302] = MEM[8310] + MEM[15372];
assign MEM[20303] = MEM[8312] + MEM[12324];
assign MEM[20304] = MEM[8313] + MEM[10549];
assign MEM[20305] = MEM[8317] + MEM[12272];
assign MEM[20306] = MEM[8318] + MEM[9016];
assign MEM[20307] = MEM[8320] + MEM[14207];
assign MEM[20308] = MEM[8321] + MEM[12505];
assign MEM[20309] = MEM[8322] + MEM[10156];
assign MEM[20310] = MEM[8323] + MEM[14081];
assign MEM[20311] = MEM[8329] + MEM[12877];
assign MEM[20312] = MEM[8330] + MEM[9255];
assign MEM[20313] = MEM[8331] + MEM[13144];
assign MEM[20314] = MEM[8336] + MEM[12573];
assign MEM[20315] = MEM[8337] + MEM[13834];
assign MEM[20316] = MEM[8338] + MEM[12900];
assign MEM[20317] = MEM[8346] + MEM[10187];
assign MEM[20318] = MEM[8347] + MEM[14341];
assign MEM[20319] = MEM[8351] + MEM[12149];
assign MEM[20320] = MEM[8352] + MEM[10070];
assign MEM[20321] = MEM[8353] + MEM[10959];
assign MEM[20322] = MEM[8354] + MEM[11426];
assign MEM[20323] = MEM[8355] + MEM[13457];
assign MEM[20324] = MEM[8356] + MEM[8492];
assign MEM[20325] = MEM[8358] + MEM[13508];
assign MEM[20326] = MEM[8360] + MEM[10917];
assign MEM[20327] = MEM[8361] + MEM[12692];
assign MEM[20328] = MEM[8365] + MEM[9142];
assign MEM[20329] = MEM[8366] + MEM[13703];
assign MEM[20330] = MEM[8383] + MEM[12941];
assign MEM[20331] = MEM[8389] + MEM[10452];
assign MEM[20332] = MEM[8394] + MEM[16267];
assign MEM[20333] = MEM[8395] + MEM[9530];
assign MEM[20334] = MEM[8398] + MEM[8817];
assign MEM[20335] = MEM[8399] + MEM[8993];
assign MEM[20336] = MEM[8400] + MEM[13317];
assign MEM[20337] = MEM[8403] + MEM[11133];
assign MEM[20338] = MEM[8404] + MEM[12561];
assign MEM[20339] = MEM[8407] + MEM[10639];
assign MEM[20340] = MEM[8410] + MEM[12679];
assign MEM[20341] = MEM[8415] + MEM[15434];
assign MEM[20342] = MEM[8417] + MEM[15859];
assign MEM[20343] = MEM[8427] + MEM[14055];
assign MEM[20344] = MEM[8428] + MEM[11523];
assign MEM[20345] = MEM[8432] + MEM[11540];
assign MEM[20346] = MEM[8434] + MEM[10226];
assign MEM[20347] = MEM[8435] + MEM[16906];
assign MEM[20348] = MEM[8436] + MEM[10911];
assign MEM[20349] = MEM[8438] + MEM[14255];
assign MEM[20350] = MEM[8440] + MEM[9131];
assign MEM[20351] = MEM[8441] + MEM[13305];
assign MEM[20352] = MEM[8443] + MEM[16949];
assign MEM[20353] = MEM[8444] + MEM[8498];
assign MEM[20354] = MEM[8445] + MEM[17086];
assign MEM[20355] = MEM[8446] + MEM[8914];
assign MEM[20356] = MEM[8454] + MEM[8518];
assign MEM[20357] = MEM[8459] + MEM[11088];
assign MEM[20358] = MEM[8460] + MEM[14827];
assign MEM[20359] = MEM[8463] + MEM[9032];
assign MEM[20360] = MEM[8468] + MEM[13976];
assign MEM[20361] = MEM[8471] + MEM[10528];
assign MEM[20362] = MEM[8475] + MEM[17418];
assign MEM[20363] = MEM[8477] + MEM[9296];
assign MEM[20364] = MEM[8478] + MEM[10092];
assign MEM[20365] = MEM[8480] + MEM[11096];
assign MEM[20366] = MEM[8481] + MEM[11895];
assign MEM[20367] = MEM[8488] + MEM[12956];
assign MEM[20368] = MEM[8491] + MEM[11999];
assign MEM[20369] = MEM[8494] + MEM[8511];
assign MEM[20370] = MEM[8495] + MEM[13780];
assign MEM[20371] = MEM[8496] + MEM[9927];
assign MEM[20372] = MEM[8500] + MEM[9816];
assign MEM[20373] = MEM[8501] + MEM[9420];
assign MEM[20374] = MEM[8503] + MEM[10203];
assign MEM[20375] = MEM[8505] + MEM[16027];
assign MEM[20376] = MEM[8506] + MEM[14191];
assign MEM[20377] = MEM[8509] + MEM[13507];
assign MEM[20378] = MEM[8515] + MEM[12535];
assign MEM[20379] = MEM[8516] + MEM[8724];
assign MEM[20380] = MEM[8519] + MEM[9603];
assign MEM[20381] = MEM[8521] + MEM[14086];
assign MEM[20382] = MEM[8522] + MEM[15180];
assign MEM[20383] = MEM[8524] + MEM[8553];
assign MEM[20384] = MEM[8528] + MEM[8917];
assign MEM[20385] = MEM[8530] + MEM[11521];
assign MEM[20386] = MEM[8531] + MEM[14889];
assign MEM[20387] = MEM[8532] + MEM[13239];
assign MEM[20388] = MEM[8538] + MEM[12156];
assign MEM[20389] = MEM[8541] + MEM[8642];
assign MEM[20390] = MEM[8542] + MEM[12810];
assign MEM[20391] = MEM[8543] + MEM[11481];
assign MEM[20392] = MEM[8544] + MEM[12559];
assign MEM[20393] = MEM[8546] + MEM[13821];
assign MEM[20394] = MEM[8549] + MEM[15156];
assign MEM[20395] = MEM[8550] + MEM[14123];
assign MEM[20396] = MEM[8555] + MEM[13036];
assign MEM[20397] = MEM[8556] + MEM[8989];
assign MEM[20398] = MEM[8561] + MEM[11361];
assign MEM[20399] = MEM[8562] + MEM[9344];
assign MEM[20400] = MEM[8567] + MEM[14672];
assign MEM[20401] = MEM[8573] + MEM[13742];
assign MEM[20402] = MEM[8575] + MEM[11204];
assign MEM[20403] = MEM[8580] + MEM[12498];
assign MEM[20404] = MEM[8581] + MEM[11041];
assign MEM[20405] = MEM[8582] + MEM[14679];
assign MEM[20406] = MEM[8583] + MEM[14576];
assign MEM[20407] = MEM[8585] + MEM[15126];
assign MEM[20408] = MEM[8587] + MEM[10254];
assign MEM[20409] = MEM[8591] + MEM[9417];
assign MEM[20410] = MEM[8596] + MEM[11349];
assign MEM[20411] = MEM[8601] + MEM[12236];
assign MEM[20412] = MEM[8604] + MEM[4786];
assign MEM[20413] = MEM[8606] + MEM[14903];
assign MEM[20414] = MEM[8607] + MEM[11256];
assign MEM[20415] = MEM[8609] + MEM[9451];
assign MEM[20416] = MEM[8618] + MEM[12117];
assign MEM[20417] = MEM[8638] + MEM[12629];
assign MEM[20418] = MEM[8644] + MEM[15344];
assign MEM[20419] = MEM[8645] + MEM[14572];
assign MEM[20420] = MEM[8652] + MEM[8718];
assign MEM[20421] = MEM[8657] + MEM[12474];
assign MEM[20422] = MEM[8661] + MEM[12386];
assign MEM[20423] = MEM[8662] + MEM[13936];
assign MEM[20424] = MEM[8663] + MEM[12347];
assign MEM[20425] = MEM[8664] + MEM[13409];
assign MEM[20426] = MEM[8665] + MEM[9037];
assign MEM[20427] = MEM[8666] + MEM[8536];
assign MEM[20428] = MEM[8670] + MEM[13895];
assign MEM[20429] = MEM[8683] + MEM[15243];
assign MEM[20430] = MEM[8687] + MEM[13377];
assign MEM[20431] = MEM[8688] + MEM[8788];
assign MEM[20432] = MEM[8690] + MEM[9866];
assign MEM[20433] = MEM[8693] + MEM[9236];
assign MEM[20434] = MEM[8694] + MEM[10654];
assign MEM[20435] = MEM[8695] + MEM[10824];
assign MEM[20436] = MEM[8696] + MEM[16660];
assign MEM[20437] = MEM[8697] + MEM[16081];
assign MEM[20438] = MEM[8698] + MEM[11062];
assign MEM[20439] = MEM[8699] + MEM[14633];
assign MEM[20440] = MEM[8704] + MEM[13014];
assign MEM[20441] = MEM[8707] + MEM[12900];
assign MEM[20442] = MEM[8708] + MEM[12907];
assign MEM[20443] = MEM[8714] + MEM[11070];
assign MEM[20444] = MEM[8719] + MEM[13333];
assign MEM[20445] = MEM[8721] + MEM[12060];
assign MEM[20446] = MEM[8725] + MEM[13571];
assign MEM[20447] = MEM[8726] + MEM[14742];
assign MEM[20448] = MEM[8727] + MEM[10835];
assign MEM[20449] = MEM[8729] + MEM[12776];
assign MEM[20450] = MEM[8730] + MEM[10712];
assign MEM[20451] = MEM[8731] + MEM[14571];
assign MEM[20452] = MEM[8732] + MEM[13252];
assign MEM[20453] = MEM[8738] + MEM[9127];
assign MEM[20454] = MEM[8740] + MEM[19656];
assign MEM[20455] = MEM[8745] + MEM[12138];
assign MEM[20456] = MEM[8749] + MEM[9564];
assign MEM[20457] = MEM[8750] + MEM[10026];
assign MEM[20458] = MEM[8761] + MEM[9996];
assign MEM[20459] = MEM[8764] + MEM[14565];
assign MEM[20460] = MEM[8768] + MEM[8922];
assign MEM[20461] = MEM[8771] + MEM[12183];
assign MEM[20462] = MEM[8773] + MEM[13323];
assign MEM[20463] = MEM[8777] + MEM[16331];
assign MEM[20464] = MEM[8780] + MEM[12620];
assign MEM[20465] = MEM[8781] + MEM[11547];
assign MEM[20466] = MEM[8783] + MEM[10895];
assign MEM[20467] = MEM[8784] + MEM[14548];
assign MEM[20468] = MEM[8786] + MEM[9267];
assign MEM[20469] = MEM[8787] + MEM[13005];
assign MEM[20470] = MEM[8792] + MEM[16771];
assign MEM[20471] = MEM[8796] + MEM[13513];
assign MEM[20472] = MEM[8799] + MEM[9116];
assign MEM[20473] = MEM[8800] + MEM[13570];
assign MEM[20474] = MEM[8801] + MEM[9017];
assign MEM[20475] = MEM[8803] + MEM[12399];
assign MEM[20476] = MEM[8804] + MEM[12073];
assign MEM[20477] = MEM[8805] + MEM[17355];
assign MEM[20478] = MEM[8816] + MEM[13168];
assign MEM[20479] = MEM[8823] + MEM[12276];
assign MEM[20480] = MEM[8824] + MEM[9456];
assign MEM[20481] = MEM[8827] + MEM[9067];
assign MEM[20482] = MEM[8828] + MEM[9184];
assign MEM[20483] = MEM[8831] + MEM[10449];
assign MEM[20484] = MEM[8834] + MEM[9908];
assign MEM[20485] = MEM[8836] + MEM[15565];
assign MEM[20486] = MEM[8837] + MEM[13555];
assign MEM[20487] = MEM[8839] + MEM[9088];
assign MEM[20488] = MEM[8841] + MEM[13511];
assign MEM[20489] = MEM[8842] + MEM[11084];
assign MEM[20490] = MEM[8845] + MEM[9061];
assign MEM[20491] = MEM[8851] + MEM[12832];
assign MEM[20492] = MEM[8857] + MEM[12327];
assign MEM[20493] = MEM[8861] + MEM[11170];
assign MEM[20494] = MEM[8862] + MEM[9950];
assign MEM[20495] = MEM[8863] + MEM[12302];
assign MEM[20496] = MEM[8865] + MEM[14645];
assign MEM[20497] = MEM[8870] + MEM[12762];
assign MEM[20498] = MEM[8875] + MEM[9422];
assign MEM[20499] = MEM[8878] + MEM[12942];
assign MEM[20500] = MEM[8883] + MEM[12017];
assign MEM[20501] = MEM[8889] + MEM[13499];
assign MEM[20502] = MEM[8891] + MEM[10728];
assign MEM[20503] = MEM[8897] + MEM[9662];
assign MEM[20504] = MEM[8907] + MEM[12898];
assign MEM[20505] = MEM[8910] + MEM[10933];
assign MEM[20506] = MEM[8919] + MEM[10717];
assign MEM[20507] = MEM[8920] + MEM[13391];
assign MEM[20508] = MEM[8923] + MEM[12153];
assign MEM[20509] = MEM[8931] + MEM[9241];
assign MEM[20510] = MEM[8934] + MEM[9674];
assign MEM[20511] = MEM[8937] + MEM[11274];
assign MEM[20512] = MEM[8938] + MEM[15012];
assign MEM[20513] = MEM[8939] + MEM[11278];
assign MEM[20514] = MEM[8941] + MEM[8962];
assign MEM[20515] = MEM[8944] + MEM[12720];
assign MEM[20516] = MEM[8948] + MEM[11783];
assign MEM[20517] = MEM[8949] + MEM[10178];
assign MEM[20518] = MEM[8951] + MEM[13365];
assign MEM[20519] = MEM[8963] + MEM[13781];
assign MEM[20520] = MEM[8968] + MEM[13077];
assign MEM[20521] = MEM[8970] + MEM[10173];
assign MEM[20522] = MEM[8972] + MEM[18122];
assign MEM[20523] = MEM[8974] + MEM[13672];
assign MEM[20524] = MEM[8975] + MEM[11346];
assign MEM[20525] = MEM[8976] + MEM[12939];
assign MEM[20526] = MEM[8978] + MEM[12442];
assign MEM[20527] = MEM[8979] + MEM[11330];
assign MEM[20528] = MEM[8981] + MEM[12139];
assign MEM[20529] = MEM[8983] + MEM[17734];
assign MEM[20530] = MEM[8986] + MEM[12196];
assign MEM[20531] = MEM[8990] + MEM[11462];
assign MEM[20532] = MEM[8997] + MEM[14939];
assign MEM[20533] = MEM[8999] + MEM[11870];
assign MEM[20534] = MEM[9002] + MEM[10161];
assign MEM[20535] = MEM[9007] + MEM[9780];
assign MEM[20536] = MEM[9009] + MEM[10125];
assign MEM[20537] = MEM[9010] + MEM[15172];
assign MEM[20538] = MEM[9011] + MEM[10761];
assign MEM[20539] = MEM[9012] + MEM[9421];
assign MEM[20540] = MEM[9013] + MEM[10076];
assign MEM[20541] = MEM[9014] + MEM[12013];
assign MEM[20542] = MEM[9018] + MEM[14488];
assign MEM[20543] = MEM[9019] + MEM[14505];
assign MEM[20544] = MEM[9020] + MEM[14157];
assign MEM[20545] = MEM[9021] + MEM[11255];
assign MEM[20546] = MEM[9024] + MEM[9828];
assign MEM[20547] = MEM[9025] + MEM[12179];
assign MEM[20548] = MEM[9026] + MEM[10578];
assign MEM[20549] = MEM[9030] + MEM[12152];
assign MEM[20550] = MEM[9031] + MEM[12366];
assign MEM[20551] = MEM[9036] + MEM[12646];
assign MEM[20552] = MEM[9038] + MEM[9122];
assign MEM[20553] = MEM[9041] + MEM[9069];
assign MEM[20554] = MEM[9042] + MEM[10861];
assign MEM[20555] = MEM[9043] + MEM[10397];
assign MEM[20556] = MEM[9044] + MEM[14238];
assign MEM[20557] = MEM[9046] + MEM[10936];
assign MEM[20558] = MEM[9051] + MEM[9229];
assign MEM[20559] = MEM[9059] + MEM[11155];
assign MEM[20560] = MEM[9060] + MEM[18241];
assign MEM[20561] = MEM[9065] + MEM[11221];
assign MEM[20562] = MEM[9070] + MEM[12488];
assign MEM[20563] = MEM[9071] + MEM[12368];
assign MEM[20564] = MEM[9073] + MEM[13218];
assign MEM[20565] = MEM[9075] + MEM[11008];
assign MEM[20566] = MEM[9076] + MEM[13321];
assign MEM[20567] = MEM[9079] + MEM[12816];
assign MEM[20568] = MEM[9082] + MEM[12828];
assign MEM[20569] = MEM[9085] + MEM[10923];
assign MEM[20570] = MEM[9087] + MEM[11173];
assign MEM[20571] = MEM[9089] + MEM[12200];
assign MEM[20572] = MEM[9090] + MEM[12631];
assign MEM[20573] = MEM[9091] + MEM[19645];
assign MEM[20574] = MEM[9092] + MEM[12577];
assign MEM[20575] = MEM[9094] + MEM[9762];
assign MEM[20576] = MEM[9095] + MEM[9381];
assign MEM[20577] = MEM[9096] + MEM[13643];
assign MEM[20578] = MEM[9099] + MEM[12903];
assign MEM[20579] = MEM[9105] + MEM[17311];
assign MEM[20580] = MEM[9107] + MEM[13245];
assign MEM[20581] = MEM[9109] + MEM[12884];
assign MEM[20582] = MEM[9111] + MEM[13671];
assign MEM[20583] = MEM[9113] + MEM[9819];
assign MEM[20584] = MEM[9114] + MEM[14204];
assign MEM[20585] = MEM[9115] + MEM[13543];
assign MEM[20586] = MEM[9117] + MEM[14533];
assign MEM[20587] = MEM[9118] + MEM[13542];
assign MEM[20588] = MEM[9120] + MEM[9494];
assign MEM[20589] = MEM[9124] + MEM[12586];
assign MEM[20590] = MEM[9126] + MEM[14756];
assign MEM[20591] = MEM[9129] + MEM[12082];
assign MEM[20592] = MEM[9132] + MEM[12129];
assign MEM[20593] = MEM[9136] + MEM[9725];
assign MEM[20594] = MEM[9140] + MEM[14646];
assign MEM[20595] = MEM[9143] + MEM[13920];
assign MEM[20596] = MEM[9144] + MEM[12100];
assign MEM[20597] = MEM[9146] + MEM[11105];
assign MEM[20598] = MEM[9150] + MEM[9211];
assign MEM[20599] = MEM[9152] + MEM[11667];
assign MEM[20600] = MEM[9153] + MEM[11061];
assign MEM[20601] = MEM[9155] + MEM[12604];
assign MEM[20602] = MEM[9158] + MEM[14553];
assign MEM[20603] = MEM[9159] + MEM[12344];
assign MEM[20604] = MEM[9161] + MEM[13289];
assign MEM[20605] = MEM[9167] + MEM[11280];
assign MEM[20606] = MEM[9168] + MEM[14110];
assign MEM[20607] = MEM[9169] + MEM[9569];
assign MEM[20608] = MEM[9170] + MEM[13946];
assign MEM[20609] = MEM[9171] + MEM[12675];
assign MEM[20610] = MEM[9172] + MEM[13774];
assign MEM[20611] = MEM[9173] + MEM[10973];
assign MEM[20612] = MEM[9177] + MEM[12006];
assign MEM[20613] = MEM[9178] + MEM[13233];
assign MEM[20614] = MEM[9179] + MEM[11318];
assign MEM[20615] = MEM[9181] + MEM[10066];
assign MEM[20616] = MEM[9186] + MEM[10997];
assign MEM[20617] = MEM[9189] + MEM[14948];
assign MEM[20618] = MEM[9190] + MEM[13606];
assign MEM[20619] = MEM[9191] + MEM[9362];
assign MEM[20620] = MEM[9194] + MEM[11177];
assign MEM[20621] = MEM[9195] + MEM[10211];
assign MEM[20622] = MEM[9197] + MEM[13436];
assign MEM[20623] = MEM[9199] + MEM[9526];
assign MEM[20624] = MEM[9200] + MEM[9214];
assign MEM[20625] = MEM[9202] + MEM[14149];
assign MEM[20626] = MEM[9215] + MEM[9846];
assign MEM[20627] = MEM[9216] + MEM[11120];
assign MEM[20628] = MEM[9217] + MEM[14051];
assign MEM[20629] = MEM[9220] + MEM[15123];
assign MEM[20630] = MEM[9221] + MEM[14899];
assign MEM[20631] = MEM[9223] + MEM[4854];
assign MEM[20632] = MEM[9224] + MEM[9463];
assign MEM[20633] = MEM[9228] + MEM[9716];
assign MEM[20634] = MEM[9232] + MEM[14836];
assign MEM[20635] = MEM[9237] + MEM[17010];
assign MEM[20636] = MEM[9238] + MEM[14617];
assign MEM[20637] = MEM[9239] + MEM[14589];
assign MEM[20638] = MEM[9246] + MEM[11711];
assign MEM[20639] = MEM[9247] + MEM[15106];
assign MEM[20640] = MEM[9250] + MEM[13509];
assign MEM[20641] = MEM[9251] + MEM[12473];
assign MEM[20642] = MEM[9252] + MEM[11902];
assign MEM[20643] = MEM[9253] + MEM[12932];
assign MEM[20644] = MEM[9256] + MEM[9489];
assign MEM[20645] = MEM[9257] + MEM[13184];
assign MEM[20646] = MEM[9260] + MEM[10948];
assign MEM[20647] = MEM[9261] + MEM[10438];
assign MEM[20648] = MEM[9262] + MEM[12133];
assign MEM[20649] = MEM[9264] + MEM[12863];
assign MEM[20650] = MEM[9266] + MEM[10601];
assign MEM[20651] = MEM[9269] + MEM[17155];
assign MEM[20652] = MEM[9271] + MEM[9774];
assign MEM[20653] = MEM[9274] + MEM[12915];
assign MEM[20654] = MEM[9280] + MEM[13080];
assign MEM[20655] = MEM[9281] + MEM[10214];
assign MEM[20656] = MEM[9284] + MEM[14173];
assign MEM[20657] = MEM[9285] + MEM[12300];
assign MEM[20658] = MEM[9286] + MEM[14045];
assign MEM[20659] = MEM[9292] + MEM[17139];
assign MEM[20660] = MEM[9293] + MEM[11716];
assign MEM[20661] = MEM[9295] + MEM[13368];
assign MEM[20662] = MEM[9297] + MEM[13170];
assign MEM[20663] = MEM[9298] + MEM[11869];
assign MEM[20664] = MEM[9300] + MEM[10108];
assign MEM[20665] = MEM[9302] + MEM[11377];
assign MEM[20666] = MEM[9305] + MEM[13414];
assign MEM[20667] = MEM[9306] + MEM[16826];
assign MEM[20668] = MEM[9307] + MEM[11130];
assign MEM[20669] = MEM[9309] + MEM[16492];
assign MEM[20670] = MEM[9314] + MEM[11179];
assign MEM[20671] = MEM[9316] + MEM[13647];
assign MEM[20672] = MEM[9318] + MEM[9804];
assign MEM[20673] = MEM[9320] + MEM[9797];
assign MEM[20674] = MEM[9322] + MEM[12796];
assign MEM[20675] = MEM[9324] + MEM[12598];
assign MEM[20676] = MEM[9329] + MEM[14369];
assign MEM[20677] = MEM[9333] + MEM[12838];
assign MEM[20678] = MEM[9334] + MEM[13854];
assign MEM[20679] = MEM[9335] + MEM[13437];
assign MEM[20680] = MEM[9336] + MEM[13679];
assign MEM[20681] = MEM[9338] + MEM[12704];
assign MEM[20682] = MEM[9340] + MEM[13471];
assign MEM[20683] = MEM[9348] + MEM[12969];
assign MEM[20684] = MEM[9349] + MEM[11350];
assign MEM[20685] = MEM[9352] + MEM[13793];
assign MEM[20686] = MEM[9353] + MEM[14787];
assign MEM[20687] = MEM[9356] + MEM[10889];
assign MEM[20688] = MEM[9358] + MEM[12536];
assign MEM[20689] = MEM[9360] + MEM[12757];
assign MEM[20690] = MEM[9364] + MEM[9759];
assign MEM[20691] = MEM[9366] + MEM[12906];
assign MEM[20692] = MEM[9368] + MEM[12261];
assign MEM[20693] = MEM[9370] + MEM[11152];
assign MEM[20694] = MEM[9372] + MEM[12916];
assign MEM[20695] = MEM[9374] + MEM[10818];
assign MEM[20696] = MEM[9377] + MEM[15921];
assign MEM[20697] = MEM[9378] + MEM[10708];
assign MEM[20698] = MEM[9384] + MEM[11031];
assign MEM[20699] = MEM[9386] + MEM[9392];
assign MEM[20700] = MEM[9389] + MEM[14108];
assign MEM[20701] = MEM[9390] + MEM[11037];
assign MEM[20702] = MEM[9391] + MEM[13068];
assign MEM[20703] = MEM[9393] + MEM[12349];
assign MEM[20704] = MEM[9395] + MEM[15950];
assign MEM[20705] = MEM[9400] + MEM[10993];
assign MEM[20706] = MEM[9404] + MEM[12656];
assign MEM[20707] = MEM[9405] + MEM[10687];
assign MEM[20708] = MEM[9408] + MEM[19984];
assign MEM[20709] = MEM[9410] + MEM[13304];
assign MEM[20710] = MEM[9412] + MEM[13146];
assign MEM[20711] = MEM[9414] + MEM[12020];
assign MEM[20712] = MEM[9418] + MEM[12146];
assign MEM[20713] = MEM[9424] + MEM[12718];
assign MEM[20714] = MEM[9425] + MEM[9681];
assign MEM[20715] = MEM[9427] + MEM[13551];
assign MEM[20716] = MEM[9428] + MEM[11187];
assign MEM[20717] = MEM[9429] + MEM[14755];
assign MEM[20718] = MEM[9431] + MEM[15091];
assign MEM[20719] = MEM[9433] + MEM[11429];
assign MEM[20720] = MEM[9434] + MEM[9510];
assign MEM[20721] = MEM[9436] + MEM[12558];
assign MEM[20722] = MEM[9437] + MEM[15296];
assign MEM[20723] = MEM[9439] + MEM[10017];
assign MEM[20724] = MEM[9441] + MEM[9997];
assign MEM[20725] = MEM[9443] + MEM[13288];
assign MEM[20726] = MEM[9444] + MEM[9642];
assign MEM[20727] = MEM[9445] + MEM[11446];
assign MEM[20728] = MEM[9446] + MEM[12143];
assign MEM[20729] = MEM[9452] + MEM[13227];
assign MEM[20730] = MEM[9457] + MEM[14744];
assign MEM[20731] = MEM[9461] + MEM[13419];
assign MEM[20732] = MEM[9467] + MEM[13094];
assign MEM[20733] = MEM[9469] + MEM[13567];
assign MEM[20734] = MEM[9470] + MEM[14723];
assign MEM[20735] = MEM[9474] + MEM[10461];
assign MEM[20736] = MEM[9477] + MEM[14427];
assign MEM[20737] = MEM[9478] + MEM[9517];
assign MEM[20738] = MEM[9482] + MEM[9932];
assign MEM[20739] = MEM[9485] + MEM[9742];
assign MEM[20740] = MEM[9490] + MEM[12777];
assign MEM[20741] = MEM[9496] + MEM[15420];
assign MEM[20742] = MEM[9498] + MEM[14034];
assign MEM[20743] = MEM[9502] + MEM[9528];
assign MEM[20744] = MEM[9504] + MEM[12418];
assign MEM[20745] = MEM[9509] + MEM[10691];
assign MEM[20746] = MEM[9511] + MEM[13673];
assign MEM[20747] = MEM[9520] + MEM[13641];
assign MEM[20748] = MEM[9523] + MEM[13370];
assign MEM[20749] = MEM[9525] + MEM[12088];
assign MEM[20750] = MEM[9529] + MEM[13206];
assign MEM[20751] = MEM[9532] + MEM[10469];
assign MEM[20752] = MEM[9538] + MEM[13782];
assign MEM[20753] = MEM[9539] + MEM[17327];
assign MEM[20754] = MEM[9541] + MEM[9679];
assign MEM[20755] = MEM[9546] + MEM[14057];
assign MEM[20756] = MEM[9549] + MEM[13985];
assign MEM[20757] = MEM[9550] + MEM[15286];
assign MEM[20758] = MEM[9553] + MEM[12355];
assign MEM[20759] = MEM[9554] + MEM[14670];
assign MEM[20760] = MEM[9557] + MEM[10755];
assign MEM[20761] = MEM[9558] + MEM[10363];
assign MEM[20762] = MEM[9559] + MEM[13721];
assign MEM[20763] = MEM[9560] + MEM[14577];
assign MEM[20764] = MEM[9562] + MEM[12808];
assign MEM[20765] = MEM[9563] + MEM[10883];
assign MEM[20766] = MEM[9566] + MEM[14094];
assign MEM[20767] = MEM[9567] + MEM[13867];
assign MEM[20768] = MEM[9570] + MEM[13250];
assign MEM[20769] = MEM[9571] + MEM[11918];
assign MEM[20770] = MEM[9572] + MEM[13790];
assign MEM[20771] = MEM[9577] + MEM[12861];
assign MEM[20772] = MEM[9578] + MEM[13657];
assign MEM[20773] = MEM[9579] + MEM[10234];
assign MEM[20774] = MEM[9580] + MEM[14350];
assign MEM[20775] = MEM[9581] + MEM[11014];
assign MEM[20776] = MEM[9583] + MEM[12118];
assign MEM[20777] = MEM[9586] + MEM[17206];
assign MEM[20778] = MEM[9590] + MEM[13791];
assign MEM[20779] = MEM[9591] + MEM[9956];
assign MEM[20780] = MEM[9597] + MEM[12281];
assign MEM[20781] = MEM[9598] + MEM[13254];
assign MEM[20782] = MEM[9600] + MEM[11142];
assign MEM[20783] = MEM[9601] + MEM[15099];
assign MEM[20784] = MEM[9604] + MEM[11302];
assign MEM[20785] = MEM[9607] + MEM[12676];
assign MEM[20786] = MEM[9618] + MEM[12013];
assign MEM[20787] = MEM[9620] + MEM[12525];
assign MEM[20788] = MEM[9622] + MEM[11497];
assign MEM[20789] = MEM[9623] + MEM[13445];
assign MEM[20790] = MEM[9626] + MEM[13691];
assign MEM[20791] = MEM[9627] + MEM[13247];
assign MEM[20792] = MEM[9633] + MEM[10428];
assign MEM[20793] = MEM[9635] + MEM[15193];
assign MEM[20794] = MEM[9638] + MEM[11022];
assign MEM[20795] = MEM[9640] + MEM[13210];
assign MEM[20796] = MEM[9641] + MEM[11259];
assign MEM[20797] = MEM[9643] + MEM[13342];
assign MEM[20798] = MEM[9644] + MEM[14962];
assign MEM[20799] = MEM[9651] + MEM[16544];
assign MEM[20800] = MEM[9652] + MEM[15930];
assign MEM[20801] = MEM[9655] + MEM[19659];
assign MEM[20802] = MEM[9660] + MEM[5746];
assign MEM[20803] = MEM[9663] + MEM[12130];
assign MEM[20804] = MEM[9664] + MEM[9921];
assign MEM[20805] = MEM[9669] + MEM[10430];
assign MEM[20806] = MEM[9671] + MEM[12016];
assign MEM[20807] = MEM[9672] + MEM[14810];
assign MEM[20808] = MEM[9673] + MEM[11132];
assign MEM[20809] = MEM[9677] + MEM[11108];
assign MEM[20810] = MEM[9678] + MEM[11598];
assign MEM[20811] = MEM[9680] + MEM[12613];
assign MEM[20812] = MEM[9682] + MEM[13002];
assign MEM[20813] = MEM[9683] + MEM[13658];
assign MEM[20814] = MEM[9686] + MEM[15377];
assign MEM[20815] = MEM[9690] + MEM[14296];
assign MEM[20816] = MEM[9692] + MEM[12697];
assign MEM[20817] = MEM[9696] + MEM[9958];
assign MEM[20818] = MEM[9697] + MEM[10760];
assign MEM[20819] = MEM[9698] + MEM[11077];
assign MEM[20820] = MEM[9699] + MEM[12681];
assign MEM[20821] = MEM[9700] + MEM[13102];
assign MEM[20822] = MEM[9701] + MEM[12829];
assign MEM[20823] = MEM[9703] + MEM[12048];
assign MEM[20824] = MEM[9705] + MEM[17158];
assign MEM[20825] = MEM[9706] + MEM[7866];
assign MEM[20826] = MEM[9710] + MEM[13336];
assign MEM[20827] = MEM[9711] + MEM[13480];
assign MEM[20828] = MEM[9715] + MEM[13488];
assign MEM[20829] = MEM[9719] + MEM[16164];
assign MEM[20830] = MEM[9720] + MEM[14901];
assign MEM[20831] = MEM[9721] + MEM[11332];
assign MEM[20832] = MEM[9724] + MEM[13429];
assign MEM[20833] = MEM[9726] + MEM[13343];
assign MEM[20834] = MEM[9728] + MEM[14195];
assign MEM[20835] = MEM[9729] + MEM[13950];
assign MEM[20836] = MEM[9730] + MEM[11536];
assign MEM[20837] = MEM[9731] + MEM[13065];
assign MEM[20838] = MEM[9736] + MEM[13496];
assign MEM[20839] = MEM[9738] + MEM[13918];
assign MEM[20840] = MEM[9740] + MEM[16965];
assign MEM[20841] = MEM[9741] + MEM[16047];
assign MEM[20842] = MEM[9744] + MEM[11571];
assign MEM[20843] = MEM[9749] + MEM[11147];
assign MEM[20844] = MEM[9751] + MEM[9973];
assign MEM[20845] = MEM[9753] + MEM[16320];
assign MEM[20846] = MEM[9757] + MEM[14367];
assign MEM[20847] = MEM[9758] + MEM[13696];
assign MEM[20848] = MEM[9760] + MEM[11229];
assign MEM[20849] = MEM[9764] + MEM[14985];
assign MEM[20850] = MEM[9765] + MEM[18338];
assign MEM[20851] = MEM[9766] + MEM[12182];
assign MEM[20852] = MEM[9767] + MEM[12831];
assign MEM[20853] = MEM[9768] + MEM[13402];
assign MEM[20854] = MEM[9769] + MEM[12299];
assign MEM[20855] = MEM[9771] + MEM[9974];
assign MEM[20856] = MEM[9772] + MEM[12683];
assign MEM[20857] = MEM[9773] + MEM[12741];
assign MEM[20858] = MEM[9777] + MEM[11471];
assign MEM[20859] = MEM[9778] + MEM[12389];
assign MEM[20860] = MEM[9781] + MEM[13385];
assign MEM[20861] = MEM[9783] + MEM[15909];
assign MEM[20862] = MEM[9784] + MEM[11378];
assign MEM[20863] = MEM[9786] + MEM[11258];
assign MEM[20864] = MEM[9787] + MEM[15428];
assign MEM[20865] = MEM[9788] + MEM[15888];
assign MEM[20866] = MEM[9789] + MEM[10662];
assign MEM[20867] = MEM[9793] + MEM[12812];
assign MEM[20868] = MEM[9794] + MEM[11976];
assign MEM[20869] = MEM[9795] + MEM[10489];
assign MEM[20870] = MEM[9798] + MEM[12781];
assign MEM[20871] = MEM[9800] + MEM[12933];
assign MEM[20872] = MEM[9801] + MEM[12752];
assign MEM[20873] = MEM[9807] + MEM[14353];
assign MEM[20874] = MEM[9814] + MEM[12329];
assign MEM[20875] = MEM[9815] + MEM[12384];
assign MEM[20876] = MEM[9818] + MEM[13320];
assign MEM[20877] = MEM[9820] + MEM[15014];
assign MEM[20878] = MEM[9821] + MEM[13023];
assign MEM[20879] = MEM[9823] + MEM[11801];
assign MEM[20880] = MEM[9824] + MEM[16392];
assign MEM[20881] = MEM[9830] + MEM[14716];
assign MEM[20882] = MEM[9831] + MEM[12644];
assign MEM[20883] = MEM[9832] + MEM[11681];
assign MEM[20884] = MEM[9833] + MEM[15953];
assign MEM[20885] = MEM[9834] + MEM[12536];
assign MEM[20886] = MEM[9835] + MEM[18804];
assign MEM[20887] = MEM[9836] + MEM[9865];
assign MEM[20888] = MEM[9839] + MEM[15326];
assign MEM[20889] = MEM[9842] + MEM[10102];
assign MEM[20890] = MEM[9844] + MEM[12297];
assign MEM[20891] = MEM[9845] + MEM[11759];
assign MEM[20892] = MEM[9848] + MEM[13899];
assign MEM[20893] = MEM[9850] + MEM[13052];
assign MEM[20894] = MEM[9851] + MEM[14833];
assign MEM[20895] = MEM[9852] + MEM[11457];
assign MEM[20896] = MEM[9854] + MEM[14214];
assign MEM[20897] = MEM[9856] + MEM[14459];
assign MEM[20898] = MEM[9858] + MEM[11127];
assign MEM[20899] = MEM[9863] + MEM[13435];
assign MEM[20900] = MEM[9864] + MEM[12976];
assign MEM[20901] = MEM[9868] + MEM[13426];
assign MEM[20902] = MEM[9872] + MEM[17250];
assign MEM[20903] = MEM[9875] + MEM[15940];
assign MEM[20904] = MEM[9876] + MEM[14162];
assign MEM[20905] = MEM[9879] + MEM[14196];
assign MEM[20906] = MEM[9881] + MEM[12363];
assign MEM[20907] = MEM[9885] + MEM[17449];
assign MEM[20908] = MEM[9886] + MEM[12826];
assign MEM[20909] = MEM[9887] + MEM[13489];
assign MEM[20910] = MEM[9893] + MEM[13820];
assign MEM[20911] = MEM[9896] + MEM[15141];
assign MEM[20912] = MEM[9897] + MEM[15414];
assign MEM[20913] = MEM[9899] + MEM[12445];
assign MEM[20914] = MEM[9904] + MEM[12985];
assign MEM[20915] = MEM[9914] + MEM[13055];
assign MEM[20916] = MEM[9915] + MEM[11385];
assign MEM[20917] = MEM[9917] + MEM[14183];
assign MEM[20918] = MEM[9918] + MEM[13371];
assign MEM[20919] = MEM[9919] + MEM[11987];
assign MEM[20920] = MEM[9922] + MEM[16210];
assign MEM[20921] = MEM[9923] + MEM[17016];
assign MEM[20922] = MEM[9924] + MEM[15568];
assign MEM[20923] = MEM[9925] + MEM[15800];
assign MEM[20924] = MEM[9926] + MEM[12700];
assign MEM[20925] = MEM[9928] + MEM[13593];
assign MEM[20926] = MEM[9930] + MEM[16003];
assign MEM[20927] = MEM[9931] + MEM[11372];
assign MEM[20928] = MEM[9937] + MEM[13183];
assign MEM[20929] = MEM[9939] + MEM[11948];
assign MEM[20930] = MEM[9940] + MEM[11515];
assign MEM[20931] = MEM[9944] + MEM[12994];
assign MEM[20932] = MEM[9947] + MEM[13994];
assign MEM[20933] = MEM[9951] + MEM[12888];
assign MEM[20934] = MEM[9952] + MEM[13891];
assign MEM[20935] = MEM[9954] + MEM[12591];
assign MEM[20936] = MEM[9959] + MEM[17124];
assign MEM[20937] = MEM[9960] + MEM[14239];
assign MEM[20938] = MEM[9962] + MEM[13131];
assign MEM[20939] = MEM[9963] + MEM[16766];
assign MEM[20940] = MEM[9965] + MEM[12986];
assign MEM[20941] = MEM[9967] + MEM[10095];
assign MEM[20942] = MEM[9969] + MEM[14541];
assign MEM[20943] = MEM[9972] + MEM[13711];
assign MEM[20944] = MEM[9978] + MEM[13381];
assign MEM[20945] = MEM[9980] + MEM[11220];
assign MEM[20946] = MEM[9982] + MEM[13098];
assign MEM[20947] = MEM[9983] + MEM[13149];
assign MEM[20948] = MEM[9984] + MEM[13659];
assign MEM[20949] = MEM[9986] + MEM[12650];
assign MEM[20950] = MEM[9988] + MEM[10981];
assign MEM[20951] = MEM[9990] + MEM[14861];
assign MEM[20952] = MEM[9991] + MEM[10544];
assign MEM[20953] = MEM[9993] + MEM[14507];
assign MEM[20954] = MEM[9999] + MEM[10216];
assign MEM[20955] = MEM[10000] + MEM[15810];
assign MEM[20956] = MEM[10003] + MEM[12643];
assign MEM[20957] = MEM[10004] + MEM[11686];
assign MEM[20958] = MEM[10009] + MEM[12926];
assign MEM[20959] = MEM[10011] + MEM[13612];
assign MEM[20960] = MEM[10012] + MEM[13617];
assign MEM[20961] = MEM[10013] + MEM[12618];
assign MEM[20962] = MEM[10014] + MEM[14503];
assign MEM[20963] = MEM[10016] + MEM[13510];
assign MEM[20964] = MEM[10020] + MEM[14069];
assign MEM[20965] = MEM[10023] + MEM[13006];
assign MEM[20966] = MEM[10025] + MEM[14032];
assign MEM[20967] = MEM[10028] + MEM[10181];
assign MEM[20968] = MEM[10029] + MEM[13880];
assign MEM[20969] = MEM[10034] + MEM[14265];
assign MEM[20970] = MEM[10035] + MEM[13058];
assign MEM[20971] = MEM[10036] + MEM[13621];
assign MEM[20972] = MEM[10043] + MEM[16773];
assign MEM[20973] = MEM[10044] + MEM[16919];
assign MEM[20974] = MEM[10048] + MEM[11466];
assign MEM[20975] = MEM[10050] + MEM[13061];
assign MEM[20976] = MEM[10051] + MEM[14457];
assign MEM[20977] = MEM[10061] + MEM[13558];
assign MEM[20978] = MEM[10064] + MEM[15993];
assign MEM[20979] = MEM[10067] + MEM[17278];
assign MEM[20980] = MEM[10072] + MEM[10905];
assign MEM[20981] = MEM[10078] + MEM[14588];
assign MEM[20982] = MEM[10079] + MEM[12075];
assign MEM[20983] = MEM[10080] + MEM[13559];
assign MEM[20984] = MEM[10082] + MEM[12237];
assign MEM[20985] = MEM[10085] + MEM[13392];
assign MEM[20986] = MEM[10086] + MEM[13294];
assign MEM[20987] = MEM[10088] + MEM[14970];
assign MEM[20988] = MEM[10089] + MEM[10256];
assign MEM[20989] = MEM[10090] + MEM[16441];
assign MEM[20990] = MEM[10091] + MEM[13945];
assign MEM[20991] = MEM[10093] + MEM[14229];
assign MEM[20992] = MEM[10094] + MEM[13404];
assign MEM[20993] = MEM[10096] + MEM[16015];
assign MEM[20994] = MEM[10100] + MEM[15669];
assign MEM[20995] = MEM[10101] + MEM[14751];
assign MEM[20996] = MEM[10103] + MEM[11928];
assign MEM[20997] = MEM[10105] + MEM[10545];
assign MEM[20998] = MEM[10106] + MEM[13515];
assign MEM[20999] = MEM[10110] + MEM[14921];
assign MEM[21000] = MEM[10116] + MEM[15814];
assign MEM[21001] = MEM[10118] + MEM[11237];
assign MEM[21002] = MEM[10121] + MEM[11005];
assign MEM[21003] = MEM[10123] + MEM[15952];
assign MEM[21004] = MEM[10124] + MEM[16936];
assign MEM[21005] = MEM[10126] + MEM[11114];
assign MEM[21006] = MEM[10132] + MEM[14006];
assign MEM[21007] = MEM[10140] + MEM[14746];
assign MEM[21008] = MEM[10141] + MEM[14725];
assign MEM[21009] = MEM[10142] + MEM[14060];
assign MEM[21010] = MEM[10144] + MEM[14963];
assign MEM[21011] = MEM[10148] + MEM[15759];
assign MEM[21012] = MEM[10153] + MEM[10400];
assign MEM[21013] = MEM[10154] + MEM[13958];
assign MEM[21014] = MEM[10155] + MEM[13362];
assign MEM[21015] = MEM[10157] + MEM[12174];
assign MEM[21016] = MEM[10160] + MEM[11925];
assign MEM[21017] = MEM[10162] + MEM[15045];
assign MEM[21018] = MEM[10164] + MEM[10570];
assign MEM[21019] = MEM[10165] + MEM[13214];
assign MEM[21020] = MEM[10166] + MEM[12165];
assign MEM[21021] = MEM[10167] + MEM[11646];
assign MEM[21022] = MEM[10169] + MEM[11823];
assign MEM[21023] = MEM[10170] + MEM[10584];
assign MEM[21024] = MEM[10171] + MEM[14967];
assign MEM[21025] = MEM[10172] + MEM[16643];
assign MEM[21026] = MEM[10176] + MEM[14599];
assign MEM[21027] = MEM[10184] + MEM[12882];
assign MEM[21028] = MEM[10188] + MEM[10998];
assign MEM[21029] = MEM[10189] + MEM[14121];
assign MEM[21030] = MEM[10191] + MEM[10957];
assign MEM[21031] = MEM[10193] + MEM[13993];
assign MEM[21032] = MEM[10195] + MEM[13020];
assign MEM[21033] = MEM[10196] + MEM[12322];
assign MEM[21034] = MEM[10198] + MEM[15134];
assign MEM[21035] = MEM[10199] + MEM[13016];
assign MEM[21036] = MEM[10201] + MEM[12633];
assign MEM[21037] = MEM[10205] + MEM[12818];
assign MEM[21038] = MEM[10212] + MEM[10546];
assign MEM[21039] = MEM[10213] + MEM[13085];
assign MEM[21040] = MEM[10215] + MEM[12811];
assign MEM[21041] = MEM[10219] + MEM[12520];
assign MEM[21042] = MEM[10225] + MEM[12780];
assign MEM[21043] = MEM[10227] + MEM[12966];
assign MEM[21044] = MEM[10231] + MEM[14542];
assign MEM[21045] = MEM[10233] + MEM[19806];
assign MEM[21046] = MEM[10235] + MEM[17808];
assign MEM[21047] = MEM[10236] + MEM[16143];
assign MEM[21048] = MEM[10238] + MEM[17852];
assign MEM[21049] = MEM[10240] + MEM[14327];
assign MEM[21050] = MEM[10242] + MEM[10576];
assign MEM[21051] = MEM[10249] + MEM[9345];
assign MEM[21052] = MEM[10251] + MEM[15543];
assign MEM[21053] = MEM[10253] + MEM[14809];
assign MEM[21054] = MEM[10258] + MEM[11416];
assign MEM[21055] = MEM[10259] + MEM[13345];
assign MEM[21056] = MEM[10261] + MEM[15055];
assign MEM[21057] = MEM[10262] + MEM[12663];
assign MEM[21058] = MEM[10263] + MEM[12189];
assign MEM[21059] = MEM[10265] + MEM[14404];
assign MEM[21060] = MEM[10266] + MEM[14300];
assign MEM[21061] = MEM[10267] + MEM[14144];
assign MEM[21062] = MEM[10269] + MEM[13330];
assign MEM[21063] = MEM[10270] + MEM[10594];
assign MEM[21064] = MEM[10274] + MEM[13042];
assign MEM[21065] = MEM[10277] + MEM[11861];
assign MEM[21066] = MEM[10277] + MEM[13982];
assign MEM[21067] = MEM[10285] + MEM[11740];
assign MEM[21068] = MEM[10287] + MEM[11154];
assign MEM[21069] = MEM[10289] + MEM[14364];
assign MEM[21070] = MEM[10293] + MEM[14281];
assign MEM[21071] = MEM[10294] + MEM[11648];
assign MEM[21072] = MEM[10296] + MEM[11013];
assign MEM[21073] = MEM[10297] + MEM[13478];
assign MEM[21074] = MEM[10298] + MEM[14113];
assign MEM[21075] = MEM[10301] + MEM[14109];
assign MEM[21076] = MEM[10302] + MEM[14895];
assign MEM[21077] = MEM[10303] + MEM[13278];
assign MEM[21078] = MEM[10305] + MEM[13681];
assign MEM[21079] = MEM[10308] + MEM[15244];
assign MEM[21080] = MEM[10310] + MEM[15264];
assign MEM[21081] = MEM[10311] + MEM[15505];
assign MEM[21082] = MEM[10312] + MEM[10814];
assign MEM[21083] = MEM[10313] + MEM[12947];
assign MEM[21084] = MEM[10314] + MEM[10561];
assign MEM[21085] = MEM[10316] + MEM[15707];
assign MEM[21086] = MEM[10317] + MEM[12560];
assign MEM[21087] = MEM[10319] + MEM[14182];
assign MEM[21088] = MEM[10326] + MEM[13076];
assign MEM[21089] = MEM[10328] + MEM[13425];
assign MEM[21090] = MEM[10329] + MEM[12514];
assign MEM[21091] = MEM[10334] + MEM[12795];
assign MEM[21092] = MEM[10335] + MEM[15519];
assign MEM[21093] = MEM[10338] + MEM[17195];
assign MEM[21094] = MEM[10340] + MEM[12820];
assign MEM[21095] = MEM[10341] + MEM[10736];
assign MEM[21096] = MEM[10342] + MEM[14640];
assign MEM[21097] = MEM[10343] + MEM[12751];
assign MEM[21098] = MEM[10344] + MEM[13473];
assign MEM[21099] = MEM[10348] + MEM[11214];
assign MEM[21100] = MEM[10349] + MEM[13150];
assign MEM[21101] = MEM[10352] + MEM[11001];
assign MEM[21102] = MEM[10355] + MEM[14030];
assign MEM[21103] = MEM[10356] + MEM[14657];
assign MEM[21104] = MEM[10357] + MEM[14821];
assign MEM[21105] = MEM[10360] + MEM[12682];
assign MEM[21106] = MEM[10361] + MEM[11248];
assign MEM[21107] = MEM[10362] + MEM[15661];
assign MEM[21108] = MEM[10364] + MEM[11911];
assign MEM[21109] = MEM[10365] + MEM[18043];
assign MEM[21110] = MEM[10372] + MEM[12693];
assign MEM[21111] = MEM[10374] + MEM[10776];
assign MEM[21112] = MEM[10375] + MEM[13819];
assign MEM[21113] = MEM[10378] + MEM[15096];
assign MEM[21114] = MEM[10379] + MEM[13257];
assign MEM[21115] = MEM[10380] + MEM[11411];
assign MEM[21116] = MEM[10384] + MEM[13275];
assign MEM[21117] = MEM[10385] + MEM[14435];
assign MEM[21118] = MEM[10387] + MEM[17337];
assign MEM[21119] = MEM[10390] + MEM[15441];
assign MEM[21120] = MEM[10394] + MEM[12911];
assign MEM[21121] = MEM[10398] + MEM[13222];
assign MEM[21122] = MEM[10401] + MEM[12213];
assign MEM[21123] = MEM[10407] + MEM[17254];
assign MEM[21124] = MEM[10408] + MEM[14201];
assign MEM[21125] = MEM[10411] + MEM[15291];
assign MEM[21126] = MEM[10412] + MEM[12494];
assign MEM[21127] = MEM[10413] + MEM[15944];
assign MEM[21128] = MEM[10416] + MEM[13154];
assign MEM[21129] = MEM[10419] + MEM[15352];
assign MEM[21130] = MEM[10420] + MEM[15408];
assign MEM[21131] = MEM[10423] + MEM[14466];
assign MEM[21132] = MEM[10425] + MEM[16345];
assign MEM[21133] = MEM[10429] + MEM[14840];
assign MEM[21134] = MEM[10436] + MEM[14528];
assign MEM[21135] = MEM[10437] + MEM[14176];
assign MEM[21136] = MEM[10441] + MEM[13814];
assign MEM[21137] = MEM[10442] + MEM[11268];
assign MEM[21138] = MEM[10447] + MEM[10604];
assign MEM[21139] = MEM[10450] + MEM[16088];
assign MEM[21140] = MEM[10455] + MEM[13539];
assign MEM[21141] = MEM[10457] + MEM[11183];
assign MEM[21142] = MEM[10458] + MEM[13461];
assign MEM[21143] = MEM[10462] + MEM[12516];
assign MEM[21144] = MEM[10471] + MEM[16096];
assign MEM[21145] = MEM[10472] + MEM[14752];
assign MEM[21146] = MEM[10484] + MEM[15356];
assign MEM[21147] = MEM[10486] + MEM[15499];
assign MEM[21148] = MEM[10488] + MEM[13686];
assign MEM[21149] = MEM[10491] + MEM[16815];
assign MEM[21150] = MEM[10493] + MEM[15022];
assign MEM[21151] = MEM[10494] + MEM[14912];
assign MEM[21152] = MEM[10496] + MEM[18554];
assign MEM[21153] = MEM[10497] + MEM[14987];
assign MEM[21154] = MEM[10499] + MEM[13879];
assign MEM[21155] = MEM[10502] + MEM[10626];
assign MEM[21156] = MEM[10504] + MEM[15367];
assign MEM[21157] = MEM[10505] + MEM[14678];
assign MEM[21158] = MEM[10507] + MEM[12873];
assign MEM[21159] = MEM[10509] + MEM[11799];
assign MEM[21160] = MEM[10512] + MEM[13477];
assign MEM[21161] = MEM[10513] + MEM[12671];
assign MEM[21162] = MEM[10514] + MEM[17126];
assign MEM[21163] = MEM[10516] + MEM[16458];
assign MEM[21164] = MEM[10517] + MEM[11320];
assign MEM[21165] = MEM[10521] + MEM[20480];
assign MEM[21166] = MEM[10525] + MEM[13029];
assign MEM[21167] = MEM[10530] + MEM[14587];
assign MEM[21168] = MEM[10533] + MEM[14283];
assign MEM[21169] = MEM[10538] + MEM[15459];
assign MEM[21170] = MEM[10539] + MEM[14893];
assign MEM[21171] = MEM[10540] + MEM[12439];
assign MEM[21172] = MEM[10542] + MEM[15581];
assign MEM[21173] = MEM[10543] + MEM[14662];
assign MEM[21174] = MEM[10548] + MEM[12909];
assign MEM[21175] = MEM[10550] + MEM[13056];
assign MEM[21176] = MEM[10552] + MEM[16699];
assign MEM[21177] = MEM[10553] + MEM[17116];
assign MEM[21178] = MEM[10562] + MEM[13779];
assign MEM[21179] = MEM[10563] + MEM[15269];
assign MEM[21180] = MEM[10564] + MEM[14063];
assign MEM[21181] = MEM[10565] + MEM[15911];
assign MEM[21182] = MEM[10569] + MEM[13758];
assign MEM[21183] = MEM[10574] + MEM[16742];
assign MEM[21184] = MEM[10575] + MEM[11289];
assign MEM[21185] = MEM[10578] + MEM[11418];
assign MEM[21186] = MEM[10582] + MEM[13619];
assign MEM[21187] = MEM[10585] + MEM[13538];
assign MEM[21188] = MEM[10590] + MEM[17008];
assign MEM[21189] = MEM[10595] + MEM[16058];
assign MEM[21190] = MEM[10597] + MEM[14531];
assign MEM[21191] = MEM[10598] + MEM[18840];
assign MEM[21192] = MEM[10601] + MEM[13996];
assign MEM[21193] = MEM[10602] + MEM[14776];
assign MEM[21194] = MEM[10603] + MEM[13875];
assign MEM[21195] = MEM[10604] + MEM[11635];
assign MEM[21196] = MEM[10606] + MEM[13828];
assign MEM[21197] = MEM[10607] + MEM[13878];
assign MEM[21198] = MEM[10609] + MEM[13767];
assign MEM[21199] = MEM[10612] + MEM[14668];
assign MEM[21200] = MEM[10615] + MEM[11786];
assign MEM[21201] = MEM[10616] + MEM[12760];
assign MEM[21202] = MEM[10617] + MEM[13923];
assign MEM[21203] = MEM[10620] + MEM[12901];
assign MEM[21204] = MEM[10624] + MEM[15445];
assign MEM[21205] = MEM[10625] + MEM[13698];
assign MEM[21206] = MEM[10627] + MEM[12162];
assign MEM[21207] = MEM[10629] + MEM[14898];
assign MEM[21208] = MEM[10631] + MEM[12202];
assign MEM[21209] = MEM[10640] + MEM[10763];
assign MEM[21210] = MEM[10645] + MEM[13706];
assign MEM[21211] = MEM[10649] + MEM[15552];
assign MEM[21212] = MEM[10654] + MEM[11574];
assign MEM[21213] = MEM[10656] + MEM[12581];
assign MEM[21214] = MEM[10658] + MEM[14007];
assign MEM[21215] = MEM[10661] + MEM[11434];
assign MEM[21216] = MEM[10661] + MEM[16361];
assign MEM[21217] = MEM[10668] + MEM[16330];
assign MEM[21218] = MEM[10671] + MEM[13598];
assign MEM[21219] = MEM[10672] + MEM[11326];
assign MEM[21220] = MEM[10674] + MEM[13125];
assign MEM[21221] = MEM[10675] + MEM[14474];
assign MEM[21222] = MEM[10678] + MEM[14357];
assign MEM[21223] = MEM[10682] + MEM[14282];
assign MEM[21224] = MEM[10683] + MEM[9515];
assign MEM[21225] = MEM[10683] + MEM[15633];
assign MEM[21226] = MEM[10686] + MEM[15877];
assign MEM[21227] = MEM[10687] + MEM[15506];
assign MEM[21228] = MEM[10689] + MEM[13948];
assign MEM[21229] = MEM[10690] + MEM[15764];
assign MEM[21230] = MEM[10693] + MEM[12833];
assign MEM[21231] = MEM[10697] + MEM[14547];
assign MEM[21232] = MEM[10720] + MEM[16476];
assign MEM[21233] = MEM[10722] + MEM[14168];
assign MEM[21234] = MEM[10725] + MEM[16698];
assign MEM[21235] = MEM[10734] + MEM[14544];
assign MEM[21236] = MEM[10735] + MEM[11109];
assign MEM[21237] = MEM[10740] + MEM[13520];
assign MEM[21238] = MEM[10746] + MEM[14402];
assign MEM[21239] = MEM[10747] + MEM[17228];
assign MEM[21240] = MEM[10762] + MEM[14624];
assign MEM[21241] = MEM[10763] + MEM[14626];
assign MEM[21242] = MEM[10772] + MEM[14686];
assign MEM[21243] = MEM[10775] + MEM[14271];
assign MEM[21244] = MEM[10777] + MEM[13850];
assign MEM[21245] = MEM[10779] + MEM[16855];
assign MEM[21246] = MEM[10785] + MEM[11125];
assign MEM[21247] = MEM[10787] + MEM[12664];
assign MEM[21248] = MEM[10790] + MEM[12622];
assign MEM[21249] = MEM[10791] + MEM[16399];
assign MEM[21250] = MEM[10800] + MEM[14740];
assign MEM[21251] = MEM[10803] + MEM[11199];
assign MEM[21252] = MEM[10803] + MEM[12733];
assign MEM[21253] = MEM[10804] + MEM[16781];
assign MEM[21254] = MEM[10806] + MEM[14140];
assign MEM[21255] = MEM[10815] + MEM[10970];
assign MEM[21256] = MEM[10815] + MEM[16412];
assign MEM[21257] = MEM[10816] + MEM[16668];
assign MEM[21258] = MEM[10817] + MEM[15103];
assign MEM[21259] = MEM[10818] + MEM[15615];
assign MEM[21260] = MEM[10822] + MEM[11267];
assign MEM[21261] = MEM[10827] + MEM[13603];
assign MEM[21262] = MEM[10828] + MEM[14496];
assign MEM[21263] = MEM[10841] + MEM[13959];
assign MEM[21264] = MEM[10842] + MEM[15991];
assign MEM[21265] = MEM[10843] + MEM[9639];
assign MEM[21266] = MEM[10847] + MEM[13246];
assign MEM[21267] = MEM[10849] + MEM[10957];
assign MEM[21268] = MEM[10852] + MEM[10988];
assign MEM[21269] = MEM[10859] + MEM[14853];
assign MEM[21270] = MEM[10863] + MEM[12905];
assign MEM[21271] = MEM[10865] + MEM[12206];
assign MEM[21272] = MEM[10866] + MEM[12899];
assign MEM[21273] = MEM[10873] + MEM[13290];
assign MEM[21274] = MEM[10880] + MEM[14432];
assign MEM[21275] = MEM[10888] + MEM[11404];
assign MEM[21276] = MEM[10888] + MEM[12360];
assign MEM[21277] = MEM[10889] + MEM[14050];
assign MEM[21278] = MEM[10890] + MEM[11672];
assign MEM[21279] = MEM[10897] + MEM[11098];
assign MEM[21280] = MEM[10900] + MEM[11545];
assign MEM[21281] = MEM[10903] + MEM[11480];
assign MEM[21282] = MEM[10907] + MEM[13863];
assign MEM[21283] = MEM[10914] + MEM[12972];
assign MEM[21284] = MEM[10924] + MEM[13518];
assign MEM[21285] = MEM[10927] + MEM[11788];
assign MEM[21286] = MEM[10933] + MEM[13833];
assign MEM[21287] = MEM[10934] + MEM[13039];
assign MEM[21288] = MEM[10943] + MEM[14857];
assign MEM[21289] = MEM[10949] + MEM[19431];
assign MEM[21290] = MEM[10954] + MEM[13565];
assign MEM[21291] = MEM[10960] + MEM[14608];
assign MEM[21292] = MEM[10965] + MEM[12885];
assign MEM[21293] = MEM[10965] + MEM[14406];
assign MEM[21294] = MEM[10971] + MEM[13132];
assign MEM[21295] = MEM[10984] + MEM[13908];
assign MEM[21296] = MEM[10985] + MEM[11718];
assign MEM[21297] = MEM[10991] + MEM[13455];
assign MEM[21298] = MEM[10999] + MEM[11696];
assign MEM[21299] = MEM[11000] + MEM[17346];
assign MEM[21300] = MEM[11017] + MEM[11617];
assign MEM[21301] = MEM[11019] + MEM[15196];
assign MEM[21302] = MEM[11026] + MEM[11390];
assign MEM[21303] = MEM[11029] + MEM[12469];
assign MEM[21304] = MEM[11029] + MEM[17192];
assign MEM[21305] = MEM[11030] + MEM[11491];
assign MEM[21306] = MEM[11034] + MEM[11441];
assign MEM[21307] = MEM[11038] + MEM[14104];
assign MEM[21308] = MEM[11039] + MEM[13156];
assign MEM[21309] = MEM[11040] + MEM[12397];
assign MEM[21310] = MEM[11043] + MEM[12067];
assign MEM[21311] = MEM[11049] + MEM[12904];
assign MEM[21312] = MEM[11054] + MEM[11067];
assign MEM[21313] = MEM[11055] + MEM[11438];
assign MEM[21314] = MEM[11059] + MEM[12325];
assign MEM[21315] = MEM[11065] + MEM[14481];
assign MEM[21316] = MEM[11078] + MEM[11376];
assign MEM[21317] = MEM[11081] + MEM[14205];
assign MEM[21318] = MEM[11083] + MEM[11257];
assign MEM[21319] = MEM[11084] + MEM[19008];
assign MEM[21320] = MEM[11086] + MEM[14513];
assign MEM[21321] = MEM[11089] + MEM[18564];
assign MEM[21322] = MEM[11091] + MEM[11236];
assign MEM[21323] = MEM[11092] + MEM[11122];
assign MEM[21324] = MEM[11097] + MEM[13083];
assign MEM[21325] = MEM[11099] + MEM[11409];
assign MEM[21326] = MEM[11104] + MEM[11980];
assign MEM[21327] = MEM[11105] + MEM[14245];
assign MEM[21328] = MEM[11106] + MEM[11126];
assign MEM[21329] = MEM[11110] + MEM[11815];
assign MEM[21330] = MEM[11112] + MEM[11964];
assign MEM[21331] = MEM[11117] + MEM[14100];
assign MEM[21332] = MEM[11118] + MEM[11794];
assign MEM[21333] = MEM[11123] + MEM[12114];
assign MEM[21334] = MEM[11128] + MEM[11145];
assign MEM[21335] = MEM[11131] + MEM[15274];
assign MEM[21336] = MEM[11134] + MEM[13155];
assign MEM[21337] = MEM[11143] + MEM[13280];
assign MEM[21338] = MEM[11144] + MEM[13423];
assign MEM[21339] = MEM[11148] + MEM[12823];
assign MEM[21340] = MEM[11164] + MEM[12121];
assign MEM[21341] = MEM[11169] + MEM[12794];
assign MEM[21342] = MEM[11170] + MEM[13632];
assign MEM[21343] = MEM[11171] + MEM[11200];
assign MEM[21344] = MEM[11174] + MEM[13067];
assign MEM[21345] = MEM[11174] + MEM[14519];
assign MEM[21346] = MEM[11176] + MEM[13212];
assign MEM[21347] = MEM[11181] + MEM[14266];
assign MEM[21348] = MEM[11182] + MEM[11217];
assign MEM[21349] = MEM[11186] + MEM[11482];
assign MEM[21350] = MEM[11188] + MEM[14262];
assign MEM[21351] = MEM[11190] + MEM[11208];
assign MEM[21352] = MEM[11191] + MEM[13616];
assign MEM[21353] = MEM[11193] + MEM[11225];
assign MEM[21354] = MEM[11194] + MEM[13710];
assign MEM[21355] = MEM[11198] + MEM[12468];
assign MEM[21356] = MEM[11202] + MEM[13303];
assign MEM[21357] = MEM[11207] + MEM[12491];
assign MEM[21358] = MEM[11209] + MEM[14165];
assign MEM[21359] = MEM[11211] + MEM[14759];
assign MEM[21360] = MEM[11213] + MEM[13729];
assign MEM[21361] = MEM[11218] + MEM[11511];
assign MEM[21362] = MEM[11226] + MEM[14040];
assign MEM[21363] = MEM[11227] + MEM[13331];
assign MEM[21364] = MEM[11230] + MEM[15226];
assign MEM[21365] = MEM[11231] + MEM[14590];
assign MEM[21366] = MEM[11233] + MEM[13277];
assign MEM[21367] = MEM[11238] + MEM[11722];
assign MEM[21368] = MEM[11240] + MEM[13632];
assign MEM[21369] = MEM[11241] + MEM[15114];
assign MEM[21370] = MEM[11246] + MEM[14390];
assign MEM[21371] = MEM[11249] + MEM[12362];
assign MEM[21372] = MEM[11262] + MEM[15704];
assign MEM[21373] = MEM[11269] + MEM[13093];
assign MEM[21374] = MEM[11270] + MEM[11329];
assign MEM[21375] = MEM[11271] + MEM[12965];
assign MEM[21376] = MEM[11273] + MEM[11444];
assign MEM[21377] = MEM[11282] + MEM[11662];
assign MEM[21378] = MEM[11284] + MEM[12991];
assign MEM[21379] = MEM[11285] + MEM[13072];
assign MEM[21380] = MEM[11293] + MEM[11430];
assign MEM[21381] = MEM[11298] + MEM[14151];
assign MEM[21382] = MEM[11299] + MEM[9403];
assign MEM[21383] = MEM[11300] + MEM[12809];
assign MEM[21384] = MEM[11307] + MEM[14619];
assign MEM[21385] = MEM[11309] + MEM[11975];
assign MEM[21386] = MEM[11313] + MEM[11857];
assign MEM[21387] = MEM[11316] + MEM[12878];
assign MEM[21388] = MEM[11319] + MEM[11506];
assign MEM[21389] = MEM[11322] + MEM[13215];
assign MEM[21390] = MEM[11323] + MEM[11250];
assign MEM[21391] = MEM[11324] + MEM[13932];
assign MEM[21392] = MEM[11325] + MEM[14998];
assign MEM[21393] = MEM[11327] + MEM[13418];
assign MEM[21394] = MEM[11331] + MEM[17395];
assign MEM[21395] = MEM[11334] + MEM[14315];
assign MEM[21396] = MEM[11335] + MEM[12393];
assign MEM[21397] = MEM[11336] + MEM[12807];
assign MEM[21398] = MEM[11337] + MEM[13799];
assign MEM[21399] = MEM[11338] + MEM[16966];
assign MEM[21400] = MEM[11339] + MEM[12840];
assign MEM[21401] = MEM[11340] + MEM[14872];
assign MEM[21402] = MEM[11341] + MEM[14320];
assign MEM[21403] = MEM[11342] + MEM[12791];
assign MEM[21404] = MEM[11347] + MEM[14476];
assign MEM[21405] = MEM[11348] + MEM[15667];
assign MEM[21406] = MEM[11353] + MEM[14303];
assign MEM[21407] = MEM[11363] + MEM[14910];
assign MEM[21408] = MEM[11364] + MEM[11654];
assign MEM[21409] = MEM[11365] + MEM[12929];
assign MEM[21410] = MEM[11366] + MEM[13253];
assign MEM[21411] = MEM[11368] + MEM[13992];
assign MEM[21412] = MEM[11369] + MEM[13805];
assign MEM[21413] = MEM[11371] + MEM[13623];
assign MEM[21414] = MEM[11373] + MEM[14116];
assign MEM[21415] = MEM[11380] + MEM[13605];
assign MEM[21416] = MEM[11381] + MEM[14348];
assign MEM[21417] = MEM[11382] + MEM[13745];
assign MEM[21418] = MEM[11384] + MEM[13845];
assign MEM[21419] = MEM[11386] + MEM[13438];
assign MEM[21420] = MEM[11387] + MEM[13099];
assign MEM[21421] = MEM[11388] + MEM[15089];
assign MEM[21422] = MEM[11392] + MEM[14150];
assign MEM[21423] = MEM[11393] + MEM[11676];
assign MEM[21424] = MEM[11394] + MEM[13964];
assign MEM[21425] = MEM[11395] + MEM[14131];
assign MEM[21426] = MEM[11397] + MEM[13637];
assign MEM[21427] = MEM[11399] + MEM[14828];
assign MEM[21428] = MEM[11400] + MEM[13866];
assign MEM[21429] = MEM[11405] + MEM[13248];
assign MEM[21430] = MEM[11410] + MEM[12889];
assign MEM[21431] = MEM[11417] + MEM[12472];
assign MEM[21432] = MEM[11419] + MEM[9514];
assign MEM[21433] = MEM[11420] + MEM[13697];
assign MEM[21434] = MEM[11424] + MEM[13561];
assign MEM[21435] = MEM[11425] + MEM[13955];
assign MEM[21436] = MEM[11427] + MEM[15563];
assign MEM[21437] = MEM[11428] + MEM[10008];
assign MEM[21438] = MEM[11432] + MEM[14983];
assign MEM[21439] = MEM[11433] + MEM[11575];
assign MEM[21440] = MEM[11435] + MEM[12448];
assign MEM[21441] = MEM[11436] + MEM[13843];
assign MEM[21442] = MEM[11440] + MEM[11538];
assign MEM[21443] = MEM[11442] + MEM[13354];
assign MEM[21444] = MEM[11445] + MEM[13823];
assign MEM[21445] = MEM[11447] + MEM[12963];
assign MEM[21446] = MEM[11449] + MEM[14031];
assign MEM[21447] = MEM[11450] + MEM[15057];
assign MEM[21448] = MEM[11453] + MEM[13807];
assign MEM[21449] = MEM[11454] + MEM[12340];
assign MEM[21450] = MEM[11455] + MEM[12522];
assign MEM[21451] = MEM[11460] + MEM[14307];
assign MEM[21452] = MEM[11461] + MEM[16816];
assign MEM[21453] = MEM[11470] + MEM[13255];
assign MEM[21454] = MEM[11472] + MEM[13204];
assign MEM[21455] = MEM[11473] + MEM[12899];
assign MEM[21456] = MEM[11475] + MEM[12728];
assign MEM[21457] = MEM[11477] + MEM[14986];
assign MEM[21458] = MEM[11484] + MEM[13947];
assign MEM[21459] = MEM[11486] + MEM[14312];
assign MEM[21460] = MEM[11488] + MEM[14099];
assign MEM[21461] = MEM[11490] + MEM[12735];
assign MEM[21462] = MEM[11492] + MEM[13186];
assign MEM[21463] = MEM[11493] + MEM[13651];
assign MEM[21464] = MEM[11495] + MEM[14133];
assign MEM[21465] = MEM[11496] + MEM[11518];
assign MEM[21466] = MEM[11499] + MEM[13595];
assign MEM[21467] = MEM[11500] + MEM[13816];
assign MEM[21468] = MEM[11503] + MEM[12294];
assign MEM[21469] = MEM[11504] + MEM[13059];
assign MEM[21470] = MEM[11507] + MEM[17420];
assign MEM[21471] = MEM[11512] + MEM[13373];
assign MEM[21472] = MEM[11513] + MEM[13261];
assign MEM[21473] = MEM[11520] + MEM[14288];
assign MEM[21474] = MEM[11522] + MEM[13315];
assign MEM[21475] = MEM[11525] + MEM[13552];
assign MEM[21476] = MEM[11526] + MEM[17268];
assign MEM[21477] = MEM[11527] + MEM[15935];
assign MEM[21478] = MEM[11528] + MEM[14663];
assign MEM[21479] = MEM[11529] + MEM[13829];
assign MEM[21480] = MEM[11531] + MEM[11860];
assign MEM[21481] = MEM[11532] + MEM[17556];
assign MEM[21482] = MEM[11533] + MEM[14860];
assign MEM[21483] = MEM[11535] + MEM[19054];
assign MEM[21484] = MEM[11542] + MEM[15436];
assign MEM[21485] = MEM[11546] + MEM[13445];
assign MEM[21486] = MEM[11549] + MEM[11636];
assign MEM[21487] = MEM[11552] + MEM[13522];
assign MEM[21488] = MEM[11553] + MEM[15333];
assign MEM[21489] = MEM[11555] + MEM[16986];
assign MEM[21490] = MEM[11557] + MEM[15027];
assign MEM[21491] = MEM[11561] + MEM[14764];
assign MEM[21492] = MEM[11568] + MEM[17057];
assign MEM[21493] = MEM[11569] + MEM[15733];
assign MEM[21494] = MEM[11574] + MEM[15382];
assign MEM[21495] = MEM[11576] + MEM[14506];
assign MEM[21496] = MEM[11578] + MEM[14246];
assign MEM[21497] = MEM[11579] + MEM[14621];
assign MEM[21498] = MEM[11580] + MEM[16607];
assign MEM[21499] = MEM[11582] + MEM[17114];
assign MEM[21500] = MEM[11584] + MEM[17458];
assign MEM[21501] = MEM[11586] + MEM[12446];
assign MEM[21502] = MEM[11591] + MEM[14444];
assign MEM[21503] = MEM[11592] + MEM[12928];
assign MEM[21504] = MEM[11593] + MEM[14349];
assign MEM[21505] = MEM[11594] + MEM[13667];
assign MEM[21506] = MEM[11600] + MEM[14187];
assign MEM[21507] = MEM[11603] + MEM[18408];
assign MEM[21508] = MEM[11604] + MEM[16978];
assign MEM[21509] = MEM[11606] + MEM[13197];
assign MEM[21510] = MEM[11607] + MEM[12817];
assign MEM[21511] = MEM[11611] + MEM[12973];
assign MEM[21512] = MEM[11612] + MEM[14391];
assign MEM[21513] = MEM[11620] + MEM[14012];
assign MEM[21514] = MEM[11626] + MEM[16601];
assign MEM[21515] = MEM[11630] + MEM[14198];
assign MEM[21516] = MEM[11633] + MEM[15176];
assign MEM[21517] = MEM[11641] + MEM[13447];
assign MEM[21518] = MEM[11642] + MEM[12582];
assign MEM[21519] = MEM[11644] + MEM[13527];
assign MEM[21520] = MEM[11645] + MEM[13279];
assign MEM[21521] = MEM[11649] + MEM[15160];
assign MEM[21522] = MEM[11650] + MEM[14516];
assign MEM[21523] = MEM[11651] + MEM[16419];
assign MEM[21524] = MEM[11656] + MEM[12109];
assign MEM[21525] = MEM[11657] + MEM[14952];
assign MEM[21526] = MEM[11659] + MEM[15313];
assign MEM[21527] = MEM[11660] + MEM[14977];
assign MEM[21528] = MEM[11661] + MEM[13648];
assign MEM[21529] = MEM[11664] + MEM[17713];
assign MEM[21530] = MEM[11670] + MEM[13979];
assign MEM[21531] = MEM[11674] + MEM[16314];
assign MEM[21532] = MEM[11678] + MEM[14661];
assign MEM[21533] = MEM[11680] + MEM[14648];
assign MEM[21534] = MEM[11682] + MEM[14438];
assign MEM[21535] = MEM[11683] + MEM[21212];
assign MEM[21536] = MEM[11688] + MEM[14793];
assign MEM[21537] = MEM[11691] + MEM[15238];
assign MEM[21538] = MEM[11692] + MEM[13636];
assign MEM[21539] = MEM[11694] + MEM[17443];
assign MEM[21540] = MEM[11695] + MEM[16921];
assign MEM[21541] = MEM[11696] + MEM[12767];
assign MEM[21542] = MEM[11698] + MEM[20974];
assign MEM[21543] = MEM[11699] + MEM[12739];
assign MEM[21544] = MEM[11703] + MEM[16799];
assign MEM[21545] = MEM[11705] + MEM[14811];
assign MEM[21546] = MEM[11708] + MEM[14338];
assign MEM[21547] = MEM[11709] + MEM[12000];
assign MEM[21548] = MEM[11712] + MEM[14130];
assign MEM[21549] = MEM[11716] + MEM[14724];
assign MEM[21550] = MEM[11717] + MEM[13633];
assign MEM[21551] = MEM[11719] + MEM[15235];
assign MEM[21552] = MEM[11721] + MEM[13972];
assign MEM[21553] = MEM[11723] + MEM[14780];
assign MEM[21554] = MEM[11726] + MEM[16648];
assign MEM[21555] = MEM[11727] + MEM[12435];
assign MEM[21556] = MEM[11728] + MEM[13674];
assign MEM[21557] = MEM[11729] + MEM[13046];
assign MEM[21558] = MEM[11731] + MEM[14114];
assign MEM[21559] = MEM[11732] + MEM[15242];
assign MEM[21560] = MEM[11733] + MEM[14882];
assign MEM[21561] = MEM[11738] + MEM[15093];
assign MEM[21562] = MEM[11739] + MEM[14504];
assign MEM[21563] = MEM[11740] + MEM[14654];
assign MEM[21564] = MEM[11747] + MEM[13358];
assign MEM[21565] = MEM[11748] + MEM[15426];
assign MEM[21566] = MEM[11750] + MEM[13422];
assign MEM[21567] = MEM[11753] + MEM[16465];
assign MEM[21568] = MEM[11756] + MEM[15742];
assign MEM[21569] = MEM[11757] + MEM[13969];
assign MEM[21570] = MEM[11758] + MEM[13336];
assign MEM[21571] = MEM[11760] + MEM[13902];
assign MEM[21572] = MEM[11761] + MEM[14344];
assign MEM[21573] = MEM[11762] + MEM[13773];
assign MEM[21574] = MEM[11764] + MEM[14945];
assign MEM[21575] = MEM[11765] + MEM[17388];
assign MEM[21576] = MEM[11767] + MEM[15200];
assign MEM[21577] = MEM[11769] + MEM[12407];
assign MEM[21578] = MEM[11770] + MEM[13203];
assign MEM[21579] = MEM[11774] + MEM[16576];
assign MEM[21580] = MEM[11776] + MEM[17081];
assign MEM[21581] = MEM[11777] + MEM[14304];
assign MEM[21582] = MEM[11779] + MEM[13274];
assign MEM[21583] = MEM[11781] + MEM[19554];
assign MEM[21584] = MEM[11785] + MEM[12690];
assign MEM[21585] = MEM[11789] + MEM[13682];
assign MEM[21586] = MEM[11802] + MEM[14943];
assign MEM[21587] = MEM[11803] + MEM[15835];
assign MEM[21588] = MEM[11804] + MEM[15677];
assign MEM[21589] = MEM[11809] + MEM[15192];
assign MEM[21590] = MEM[11810] + MEM[14779];
assign MEM[21591] = MEM[11811] + MEM[12533];
assign MEM[21592] = MEM[11812] + MEM[12685];
assign MEM[21593] = MEM[11816] + MEM[15214];
assign MEM[21594] = MEM[11818] + MEM[14248];
assign MEM[21595] = MEM[11820] + MEM[16246];
assign MEM[21596] = MEM[11821] + MEM[12769];
assign MEM[21597] = MEM[11824] + MEM[13504];
assign MEM[21598] = MEM[11825] + MEM[13761];
assign MEM[21599] = MEM[11827] + MEM[14612];
assign MEM[21600] = MEM[11828] + MEM[15992];
assign MEM[21601] = MEM[11829] + MEM[15150];
assign MEM[21602] = MEM[11830] + MEM[12888];
assign MEM[21603] = MEM[11835] + MEM[14434];
assign MEM[21604] = MEM[11836] + MEM[15017];
assign MEM[21605] = MEM[11842] + MEM[12362];
assign MEM[21606] = MEM[11843] + MEM[13417];
assign MEM[21607] = MEM[11850] + MEM[15036];
assign MEM[21608] = MEM[11852] + MEM[14647];
assign MEM[21609] = MEM[11858] + MEM[15288];
assign MEM[21610] = MEM[11859] + MEM[20150];
assign MEM[21611] = MEM[11871] + MEM[12017];
assign MEM[21612] = MEM[11872] + MEM[13450];
assign MEM[21613] = MEM[11875] + MEM[15257];
assign MEM[21614] = MEM[11878] + MEM[13811];
assign MEM[21615] = MEM[11881] + MEM[9593];
assign MEM[21616] = MEM[11884] + MEM[15582];
assign MEM[21617] = MEM[11886] + MEM[16033];
assign MEM[21618] = MEM[11888] + MEM[13915];
assign MEM[21619] = MEM[11891] + MEM[15157];
assign MEM[21620] = MEM[11894] + MEM[14512];
assign MEM[21621] = MEM[11896] + MEM[15390];
assign MEM[21622] = MEM[11900] + MEM[17129];
assign MEM[21623] = MEM[11903] + MEM[19487];
assign MEM[21624] = MEM[11904] + MEM[13129];
assign MEM[21625] = MEM[11906] + MEM[14156];
assign MEM[21626] = MEM[11908] + MEM[14268];
assign MEM[21627] = MEM[11912] + MEM[14103];
assign MEM[21628] = MEM[11913] + MEM[16473];
assign MEM[21629] = MEM[11920] + MEM[13573];
assign MEM[21630] = MEM[11921] + MEM[18569];
assign MEM[21631] = MEM[11927] + MEM[16929];
assign MEM[21632] = MEM[11941] + MEM[16311];
assign MEM[21633] = MEM[11947] + MEM[15066];
assign MEM[21634] = MEM[11949] + MEM[15840];
assign MEM[21635] = MEM[11951] + MEM[18381];
assign MEM[21636] = MEM[11952] + MEM[14232];
assign MEM[21637] = MEM[11953] + MEM[15985];
assign MEM[21638] = MEM[11956] + MEM[15061];
assign MEM[21639] = MEM[11968] + MEM[14453];
assign MEM[21640] = MEM[11970] + MEM[14848];
assign MEM[21641] = MEM[11971] + MEM[14362];
assign MEM[21642] = MEM[11972] + MEM[13353];
assign MEM[21643] = MEM[11974] + MEM[12364];
assign MEM[21644] = MEM[11978] + MEM[14942];
assign MEM[21645] = MEM[11983] + MEM[17361];
assign MEM[21646] = MEM[11984] + MEM[14675];
assign MEM[21647] = MEM[11986] + MEM[16708];
assign MEM[21648] = MEM[11988] + MEM[20701];
assign MEM[21649] = MEM[11996] + MEM[15136];
assign MEM[21650] = MEM[12003] + MEM[13921];
assign MEM[21651] = MEM[12004] + MEM[13900];
assign MEM[21652] = MEM[12005] + MEM[13720];
assign MEM[21653] = MEM[12008] + MEM[17451];
assign MEM[21654] = MEM[12010] + MEM[15021];
assign MEM[21655] = MEM[12012] + MEM[14574];
assign MEM[21656] = MEM[12014] + MEM[13335];
assign MEM[21657] = MEM[12015] + MEM[15217];
assign MEM[21658] = MEM[12018] + MEM[17576];
assign MEM[21659] = MEM[12021] + MEM[15237];
assign MEM[21660] = MEM[12023] + MEM[16870];
assign MEM[21661] = MEM[12024] + MEM[14824];
assign MEM[21662] = MEM[12027] + MEM[14482];
assign MEM[21663] = MEM[12028] + MEM[20697];
assign MEM[21664] = MEM[12029] + MEM[12660];
assign MEM[21665] = MEM[12030] + MEM[15000];
assign MEM[21666] = MEM[12032] + MEM[13926];
assign MEM[21667] = MEM[12035] + MEM[14403];
assign MEM[21668] = MEM[12036] + MEM[14172];
assign MEM[21669] = MEM[12038] + MEM[16409];
assign MEM[21670] = MEM[12039] + MEM[12775];
assign MEM[21671] = MEM[12041] + MEM[16755];
assign MEM[21672] = MEM[12042] + MEM[13166];
assign MEM[21673] = MEM[12043] + MEM[14522];
assign MEM[21674] = MEM[12044] + MEM[12930];
assign MEM[21675] = MEM[12045] + MEM[12949];
assign MEM[21676] = MEM[12049] + MEM[15336];
assign MEM[21677] = MEM[12051] + MEM[17391];
assign MEM[21678] = MEM[12052] + MEM[14768];
assign MEM[21679] = MEM[12054] + MEM[14774];
assign MEM[21680] = MEM[12055] + MEM[12855];
assign MEM[21681] = MEM[12063] + MEM[15391];
assign MEM[21682] = MEM[12065] + MEM[14859];
assign MEM[21683] = MEM[12066] + MEM[12927];
assign MEM[21684] = MEM[12071] + MEM[15026];
assign MEM[21685] = MEM[12072] + MEM[12657];
assign MEM[21686] = MEM[12076] + MEM[14065];
assign MEM[21687] = MEM[12077] + MEM[14789];
assign MEM[21688] = MEM[12078] + MEM[15907];
assign MEM[21689] = MEM[12082] + MEM[17437];
assign MEM[21690] = MEM[12083] + MEM[20372];
assign MEM[21691] = MEM[12084] + MEM[9325];
assign MEM[21692] = MEM[12092] + MEM[18391];
assign MEM[21693] = MEM[12100] + MEM[19283];
assign MEM[21694] = MEM[12103] + MEM[16174];
assign MEM[21695] = MEM[12109] + MEM[14376];
assign MEM[21696] = MEM[12118] + MEM[14247];
assign MEM[21697] = MEM[12128] + MEM[12553];
assign MEM[21698] = MEM[12137] + MEM[17221];
assign MEM[21699] = MEM[12139] + MEM[14781];
assign MEM[21700] = MEM[12144] + MEM[13108];
assign MEM[21701] = MEM[12146] + MEM[15232];
assign MEM[21702] = MEM[12157] + MEM[14530];
assign MEM[21703] = MEM[12160] + MEM[13019];
assign MEM[21704] = MEM[12161] + MEM[15102];
assign MEM[21705] = MEM[12165] + MEM[17478];
assign MEM[21706] = MEM[12166] + MEM[14914];
assign MEM[21707] = MEM[12174] + MEM[12471];
assign MEM[21708] = MEM[12183] + MEM[15087];
assign MEM[21709] = MEM[12185] + MEM[13226];
assign MEM[21710] = MEM[12188] + MEM[15856];
assign MEM[21711] = MEM[12189] + MEM[16167];
assign MEM[21712] = MEM[12192] + MEM[12210];
assign MEM[21713] = MEM[12205] + MEM[14372];
assign MEM[21714] = MEM[12206] + MEM[13930];
assign MEM[21715] = MEM[12218] + MEM[15228];
assign MEM[21716] = MEM[12219] + MEM[17399];
assign MEM[21717] = MEM[12220] + MEM[14480];
assign MEM[21718] = MEM[12225] + MEM[15458];
assign MEM[21719] = MEM[12227] + MEM[18102];
assign MEM[21720] = MEM[12232] + MEM[17060];
assign MEM[21721] = MEM[12245] + MEM[16055];
assign MEM[21722] = MEM[12252] + MEM[15060];
assign MEM[21723] = MEM[12256] + MEM[14431];
assign MEM[21724] = MEM[12263] + MEM[13707];
assign MEM[21725] = MEM[12263] + MEM[17251];
assign MEM[21726] = MEM[12265] + MEM[15734];
assign MEM[21727] = MEM[12268] + MEM[14073];
assign MEM[21728] = MEM[12272] + MEM[15648];
assign MEM[21729] = MEM[12273] + MEM[13316];
assign MEM[21730] = MEM[12276] + MEM[15325];
assign MEM[21731] = MEM[12277] + MEM[16652];
assign MEM[21732] = MEM[12278] + MEM[15004];
assign MEM[21733] = MEM[12281] + MEM[13903];
assign MEM[21734] = MEM[12282] + MEM[13201];
assign MEM[21735] = MEM[12282] + MEM[13287];
assign MEM[21736] = MEM[12283] + MEM[14154];
assign MEM[21737] = MEM[12284] + MEM[15400];
assign MEM[21738] = MEM[12285] + MEM[13272];
assign MEM[21739] = MEM[12286] + MEM[17842];
assign MEM[21740] = MEM[12296] + MEM[16105];
assign MEM[21741] = MEM[12297] + MEM[16226];
assign MEM[21742] = MEM[12299] + MEM[14613];
assign MEM[21743] = MEM[12300] + MEM[15148];
assign MEM[21744] = MEM[12308] + MEM[16178];
assign MEM[21745] = MEM[12311] + MEM[13835];
assign MEM[21746] = MEM[12312] + MEM[15202];
assign MEM[21747] = MEM[12319] + MEM[13544];
assign MEM[21748] = MEM[12324] + MEM[13725];
assign MEM[21749] = MEM[12325] + MEM[14142];
assign MEM[21750] = MEM[12329] + MEM[14087];
assign MEM[21751] = MEM[12333] + MEM[15685];
assign MEM[21752] = MEM[12334] + MEM[14382];
assign MEM[21753] = MEM[12335] + MEM[17184];
assign MEM[21754] = MEM[12341] + MEM[15083];
assign MEM[21755] = MEM[12342] + MEM[13177];
assign MEM[21756] = MEM[12345] + MEM[14383];
assign MEM[21757] = MEM[12347] + MEM[17392];
assign MEM[21758] = MEM[12350] + MEM[14462];
assign MEM[21759] = MEM[12351] + MEM[15891];
assign MEM[21760] = MEM[12363] + MEM[13700];
assign MEM[21761] = MEM[12366] + MEM[15711];
assign MEM[21762] = MEM[12369] + MEM[13384];
assign MEM[21763] = MEM[12373] + MEM[14036];
assign MEM[21764] = MEM[12375] + MEM[16776];
assign MEM[21765] = MEM[12380] + MEM[13217];
assign MEM[21766] = MEM[12380] + MEM[16907];
assign MEM[21767] = MEM[12381] + MEM[17532];
assign MEM[21768] = MEM[12386] + MEM[15621];
assign MEM[21769] = MEM[12387] + MEM[14635];
assign MEM[21770] = MEM[12388] + MEM[15182];
assign MEM[21771] = MEM[12388] + MEM[18076];
assign MEM[21772] = MEM[12391] + MEM[13694];
assign MEM[21773] = MEM[12391] + MEM[13927];
assign MEM[21774] = MEM[12393] + MEM[16737];
assign MEM[21775] = MEM[12395] + MEM[12465];
assign MEM[21776] = MEM[12407] + MEM[15316];
assign MEM[21777] = MEM[12413] + MEM[16690];
assign MEM[21778] = MEM[12418] + MEM[14991];
assign MEM[21779] = MEM[12425] + MEM[15657];
assign MEM[21780] = MEM[12426] + MEM[14375];
assign MEM[21781] = MEM[12430] + MEM[13059];
assign MEM[21782] = MEM[12444] + MEM[13265];
assign MEM[21783] = MEM[12447] + MEM[15236];
assign MEM[21784] = MEM[12453] + MEM[13172];
assign MEM[21785] = MEM[12455] + MEM[14186];
assign MEM[21786] = MEM[12460] + MEM[17204];
assign MEM[21787] = MEM[12462] + MEM[13281];
assign MEM[21788] = MEM[12463] + MEM[14747];
assign MEM[21789] = MEM[12469] + MEM[15412];
assign MEM[21790] = MEM[12473] + MEM[17244];
assign MEM[21791] = MEM[12474] + MEM[16244];
assign MEM[21792] = MEM[12478] + MEM[14845];
assign MEM[21793] = MEM[12480] + MEM[14251];
assign MEM[21794] = MEM[12481] + MEM[14306];
assign MEM[21795] = MEM[12487] + MEM[14458];
assign MEM[21796] = MEM[12494] + MEM[17731];
assign MEM[21797] = MEM[12499] + MEM[13735];
assign MEM[21798] = MEM[12504] + MEM[14351];
assign MEM[21799] = MEM[12506] + MEM[13842];
assign MEM[21800] = MEM[12512] + MEM[19724];
assign MEM[21801] = MEM[12514] + MEM[16559];
assign MEM[21802] = MEM[12518] + MEM[12591];
assign MEM[21803] = MEM[12524] + MEM[16116];
assign MEM[21804] = MEM[12531] + MEM[13080];
assign MEM[21805] = MEM[12533] + MEM[20703];
assign MEM[21806] = MEM[12537] + MEM[15334];
assign MEM[21807] = MEM[12538] + MEM[12566];
assign MEM[21808] = MEM[12544] + MEM[12925];
assign MEM[21809] = MEM[12555] + MEM[13595];
assign MEM[21810] = MEM[12557] + MEM[15249];
assign MEM[21811] = MEM[12558] + MEM[14269];
assign MEM[21812] = MEM[12560] + MEM[20278];
assign MEM[21813] = MEM[12566] + MEM[13890];
assign MEM[21814] = MEM[12573] + MEM[14949];
assign MEM[21815] = MEM[12576] + MEM[15936];
assign MEM[21816] = MEM[12577] + MEM[12584];
assign MEM[21817] = MEM[12583] + MEM[15404];
assign MEM[21818] = MEM[12593] + MEM[17299];
assign MEM[21819] = MEM[12599] + MEM[15129];
assign MEM[21820] = MEM[12610] + MEM[8640];
assign MEM[21821] = MEM[12610] + MEM[15271];
assign MEM[21822] = MEM[12612] + MEM[14753];
assign MEM[21823] = MEM[12622] + MEM[14171];
assign MEM[21824] = MEM[12623] + MEM[14047];
assign MEM[21825] = MEM[12624] + MEM[14439];
assign MEM[21826] = MEM[12626] + MEM[17161];
assign MEM[21827] = MEM[12628] + MEM[12646];
assign MEM[21828] = MEM[12629] + MEM[17409];
assign MEM[21829] = MEM[12643] + MEM[18404];
assign MEM[21830] = MEM[12644] + MEM[15056];
assign MEM[21831] = MEM[12645] + MEM[14674];
assign MEM[21832] = MEM[12656] + MEM[14796];
assign MEM[21833] = MEM[12660] + MEM[15465];
assign MEM[21834] = MEM[12663] + MEM[14380];
assign MEM[21835] = MEM[12664] + MEM[15357];
assign MEM[21836] = MEM[12666] + MEM[13140];
assign MEM[21837] = MEM[12671] + MEM[14696];
assign MEM[21838] = MEM[12674] + MEM[14524];
assign MEM[21839] = MEM[12686] + MEM[14642];
assign MEM[21840] = MEM[12692] + MEM[16938];
assign MEM[21841] = MEM[12699] + MEM[12897];
assign MEM[21842] = MEM[12699] + MEM[14920];
assign MEM[21843] = MEM[12701] + MEM[13795];
assign MEM[21844] = MEM[12709] + MEM[19114];
assign MEM[21845] = MEM[12710] + MEM[13680];
assign MEM[21846] = MEM[12711] + MEM[13718];
assign MEM[21847] = MEM[12722] + MEM[15204];
assign MEM[21848] = MEM[12727] + MEM[12904];
assign MEM[21849] = MEM[12732] + MEM[13603];
assign MEM[21850] = MEM[12733] + MEM[17283];
assign MEM[21851] = MEM[12734] + MEM[15041];
assign MEM[21852] = MEM[12737] + MEM[14815];
assign MEM[21853] = MEM[12739] + MEM[14465];
assign MEM[21854] = MEM[12741] + MEM[15539];
assign MEM[21855] = MEM[12749] + MEM[15342];
assign MEM[21856] = MEM[12750] + MEM[17233];
assign MEM[21857] = MEM[12755] + MEM[13387];
assign MEM[21858] = MEM[12760] + MEM[14261];
assign MEM[21859] = MEM[12763] + MEM[14072];
assign MEM[21860] = MEM[12770] + MEM[13748];
assign MEM[21861] = MEM[12772] + MEM[19994];
assign MEM[21862] = MEM[12773] + MEM[13139];
assign MEM[21863] = MEM[12774] + MEM[17243];
assign MEM[21864] = MEM[12775] + MEM[15945];
assign MEM[21865] = MEM[12776] + MEM[14975];
assign MEM[21866] = MEM[12777] + MEM[20592];
assign MEM[21867] = MEM[12780] + MEM[15149];
assign MEM[21868] = MEM[12784] + MEM[15327];
assign MEM[21869] = MEM[12785] + MEM[16068];
assign MEM[21870] = MEM[12786] + MEM[15647];
assign MEM[21871] = MEM[12790] + MEM[14673];
assign MEM[21872] = MEM[12790] + MEM[14019];
assign MEM[21873] = MEM[12795] + MEM[16036];
assign MEM[21874] = MEM[12796] + MEM[14748];
assign MEM[21875] = MEM[12799] + MEM[13913];
assign MEM[21876] = MEM[12807] + MEM[14600];
assign MEM[21877] = MEM[12810] + MEM[14551];
assign MEM[21878] = MEM[12811] + MEM[13176];
assign MEM[21879] = MEM[12813] + MEM[13358];
assign MEM[21880] = MEM[12815] + MEM[13962];
assign MEM[21881] = MEM[12818] + MEM[15298];
assign MEM[21882] = MEM[12820] + MEM[13017];
assign MEM[21883] = MEM[12823] + MEM[14813];
assign MEM[21884] = MEM[12831] + MEM[17477];
assign MEM[21885] = MEM[12832] + MEM[14398];
assign MEM[21886] = MEM[12833] + MEM[15388];
assign MEM[21887] = MEM[12835] + MEM[15901];
assign MEM[21888] = MEM[12840] + MEM[14228];
assign MEM[21889] = MEM[12844] + MEM[14276];
assign MEM[21890] = MEM[12849] + MEM[13844];
assign MEM[21891] = MEM[12856] + MEM[14867];
assign MEM[21892] = MEM[12856] + MEM[15393];
assign MEM[21893] = MEM[12862] + MEM[15872];
assign MEM[21894] = MEM[12873] + MEM[14250];
assign MEM[21895] = MEM[12879] + MEM[13223];
assign MEM[21896] = MEM[12884] + MEM[15023];
assign MEM[21897] = MEM[12885] + MEM[17012];
assign MEM[21898] = MEM[12886] + MEM[13168];
assign MEM[21899] = MEM[12887] + MEM[13560];
assign MEM[21900] = MEM[12889] + MEM[13375];
assign MEM[21901] = MEM[12893] + MEM[17276];
assign MEM[21902] = MEM[12897] + MEM[13661];
assign MEM[21903] = MEM[12898] + MEM[14667];
assign MEM[21904] = MEM[12902] + MEM[13377];
assign MEM[21905] = MEM[12907] + MEM[14990];
assign MEM[21906] = MEM[12908] + MEM[15130];
assign MEM[21907] = MEM[12909] + MEM[19926];
assign MEM[21908] = MEM[12915] + MEM[15062];
assign MEM[21909] = MEM[12916] + MEM[13601];
assign MEM[21910] = MEM[12917] + MEM[13069];
assign MEM[21911] = MEM[12921] + MEM[13137];
assign MEM[21912] = MEM[12931] + MEM[15019];
assign MEM[21913] = MEM[12937] + MEM[14979];
assign MEM[21914] = MEM[12939] + MEM[21185];
assign MEM[21915] = MEM[12941] + MEM[15688];
assign MEM[21916] = MEM[12942] + MEM[14880];
assign MEM[21917] = MEM[12949] + MEM[16940];
assign MEM[21918] = MEM[12953] + MEM[15178];
assign MEM[21919] = MEM[12956] + MEM[14790];
assign MEM[21920] = MEM[12961] + MEM[13584];
assign MEM[21921] = MEM[12965] + MEM[14736];
assign MEM[21922] = MEM[12966] + MEM[14549];
assign MEM[21923] = MEM[12982] + MEM[13041];
assign MEM[21924] = MEM[12982] + MEM[17091];
assign MEM[21925] = MEM[12983] + MEM[13557];
assign MEM[21926] = MEM[12984] + MEM[13609];
assign MEM[21927] = MEM[12984] + MEM[15152];
assign MEM[21928] = MEM[12985] + MEM[19579];
assign MEM[21929] = MEM[12986] + MEM[15592];
assign MEM[21930] = MEM[12991] + MEM[14800];
assign MEM[21931] = MEM[12997] + MEM[14412];
assign MEM[21932] = MEM[13005] + MEM[15266];
assign MEM[21933] = MEM[13009] + MEM[18635];
assign MEM[21934] = MEM[13014] + MEM[14192];
assign MEM[21935] = MEM[13020] + MEM[15268];
assign MEM[21936] = MEM[13021] + MEM[13389];
assign MEM[21937] = MEM[13023] + MEM[13858];
assign MEM[21938] = MEM[13024] + MEM[13712];
assign MEM[21939] = MEM[13027] + MEM[14139];
assign MEM[21940] = MEM[13030] + MEM[14025];
assign MEM[21941] = MEM[13032] + MEM[14597];
assign MEM[21942] = MEM[13033] + MEM[13970];
assign MEM[21943] = MEM[13036] + MEM[14336];
assign MEM[21944] = MEM[13040] + MEM[3942];
assign MEM[21945] = MEM[13041] + MEM[13980];
assign MEM[21946] = MEM[13044] + MEM[13314];
assign MEM[21947] = MEM[13047] + MEM[9599];
assign MEM[21948] = MEM[13048] + MEM[19247];
assign MEM[21949] = MEM[13053] + MEM[13702];
assign MEM[21950] = MEM[13053] + MEM[16076];
assign MEM[21951] = MEM[13055] + MEM[19803];
assign MEM[21952] = MEM[13057] + MEM[14164];
assign MEM[21953] = MEM[13057] + MEM[15115];
assign MEM[21954] = MEM[13060] + MEM[15425];
assign MEM[21955] = MEM[13066] + MEM[14726];
assign MEM[21956] = MEM[13067] + MEM[15159];
assign MEM[21957] = MEM[13070] + MEM[13824];
assign MEM[21958] = MEM[13070] + MEM[15037];
assign MEM[21959] = MEM[13074] + MEM[13628];
assign MEM[21960] = MEM[13081] + MEM[13186];
assign MEM[21961] = MEM[13086] + MEM[17945];
assign MEM[21962] = MEM[13087] + MEM[9491];
assign MEM[21963] = MEM[13087] + MEM[15915];
assign MEM[21964] = MEM[13092] + MEM[15447];
assign MEM[21965] = MEM[13094] + MEM[15916];
assign MEM[21966] = MEM[13099] + MEM[15024];
assign MEM[21967] = MEM[13104] + MEM[13690];
assign MEM[21968] = MEM[13108] + MEM[13563];
assign MEM[21969] = MEM[13110] + MEM[13260];
assign MEM[21970] = MEM[13115] + MEM[16814];
assign MEM[21971] = MEM[13116] + MEM[14433];
assign MEM[21972] = MEM[13117] + MEM[15133];
assign MEM[21973] = MEM[13131] + MEM[13479];
assign MEM[21974] = MEM[13133] + MEM[14713];
assign MEM[21975] = MEM[13137] + MEM[16084];
assign MEM[21976] = MEM[13144] + MEM[14016];
assign MEM[21977] = MEM[13146] + MEM[15127];
assign MEM[21978] = MEM[13147] + MEM[14883];
assign MEM[21979] = MEM[13151] + MEM[15775];
assign MEM[21980] = MEM[13153] + MEM[14128];
assign MEM[21981] = MEM[13155] + MEM[15030];
assign MEM[21982] = MEM[13161] + MEM[16729];
assign MEM[21983] = MEM[13166] + MEM[13737];
assign MEM[21984] = MEM[13167] + MEM[13594];
assign MEM[21985] = MEM[13169] + MEM[14408];
assign MEM[21986] = MEM[13169] + MEM[20355];
assign MEM[21987] = MEM[13171] + MEM[19260];
assign MEM[21988] = MEM[13172] + MEM[15005];
assign MEM[21989] = MEM[13174] + MEM[14450];
assign MEM[21990] = MEM[13174] + MEM[15285];
assign MEM[21991] = MEM[13179] + MEM[15281];
assign MEM[21992] = MEM[13183] + MEM[14360];
assign MEM[21993] = MEM[13185] + MEM[13363];
assign MEM[21994] = MEM[13185] + MEM[15065];
assign MEM[21995] = MEM[13194] + MEM[15491];
assign MEM[21996] = MEM[13197] + MEM[14688];
assign MEM[21997] = MEM[13198] + MEM[14495];
assign MEM[21998] = MEM[13201] + MEM[14294];
assign MEM[21999] = MEM[13202] + MEM[18742];
assign MEM[22000] = MEM[13203] + MEM[13754];
assign MEM[22001] = MEM[13213] + MEM[14352];
assign MEM[22002] = MEM[13213] + MEM[14414];
assign MEM[22003] = MEM[13214] + MEM[15655];
assign MEM[22004] = MEM[13216] + MEM[14812];
assign MEM[22005] = MEM[13218] + MEM[17095];
assign MEM[22006] = MEM[13222] + MEM[16817];
assign MEM[22007] = MEM[13228] + MEM[13649];
assign MEM[22008] = MEM[13229] + MEM[13638];
assign MEM[22009] = MEM[13231] + MEM[13475];
assign MEM[22010] = MEM[13233] + MEM[16667];
assign MEM[22011] = MEM[13238] + MEM[13770];
assign MEM[22012] = MEM[13238] + MEM[17135];
assign MEM[22013] = MEM[13239] + MEM[15340];
assign MEM[22014] = MEM[13240] + MEM[14908];
assign MEM[22015] = MEM[13253] + MEM[15112];
assign MEM[22016] = MEM[13254] + MEM[16004];
assign MEM[22017] = MEM[13260] + MEM[13561];
assign MEM[22018] = MEM[13261] + MEM[16794];
assign MEM[22019] = MEM[13262] + MEM[13655];
assign MEM[22020] = MEM[13262] + MEM[16487];
assign MEM[22021] = MEM[13265] + MEM[16250];
assign MEM[22022] = MEM[13266] + MEM[15310];
assign MEM[22023] = MEM[13267] + MEM[13394];
assign MEM[22024] = MEM[13270] + MEM[14944];
assign MEM[22025] = MEM[13274] + MEM[13931];
assign MEM[22026] = MEM[13275] + MEM[20017];
assign MEM[22027] = MEM[13289] + MEM[16454];
assign MEM[22028] = MEM[13295] + MEM[13532];
assign MEM[22029] = MEM[13302] + MEM[13378];
assign MEM[22030] = MEM[13302] + MEM[21082];
assign MEM[22031] = MEM[13303] + MEM[18601];
assign MEM[22032] = MEM[13306] + MEM[14839];
assign MEM[22033] = MEM[13310] + MEM[13699];
assign MEM[22034] = MEM[13312] + MEM[15725];
assign MEM[22035] = MEM[13316] + MEM[13648];
assign MEM[22036] = MEM[13320] + MEM[15137];
assign MEM[22037] = MEM[13321] + MEM[15440];
assign MEM[22038] = MEM[13322] + MEM[14956];
assign MEM[22039] = MEM[13323] + MEM[14799];
assign MEM[22040] = MEM[13343] + MEM[14708];
assign MEM[22041] = MEM[13345] + MEM[17431];
assign MEM[22042] = MEM[13353] + MEM[15218];
assign MEM[22043] = MEM[13356] + MEM[21510];
assign MEM[22044] = MEM[13359] + MEM[14849];
assign MEM[22045] = MEM[13359] + MEM[14924];
assign MEM[22046] = MEM[13376] + MEM[15046];
assign MEM[22047] = MEM[13379] + MEM[14644];
assign MEM[22048] = MEM[13384] + MEM[17220];
assign MEM[22049] = MEM[13388] + MEM[13777];
assign MEM[22050] = MEM[13388] + MEM[16976];
assign MEM[22051] = MEM[13395] + MEM[20457];
assign MEM[22052] = MEM[13398] + MEM[14274];
assign MEM[22053] = MEM[13398] + MEM[15757];
assign MEM[22054] = MEM[13400] + MEM[15201];
assign MEM[22055] = MEM[13401] + MEM[14329];
assign MEM[22056] = MEM[13406] + MEM[13798];
assign MEM[22057] = MEM[13414] + MEM[15307];
assign MEM[22058] = MEM[13415] + MEM[13645];
assign MEM[22059] = MEM[13415] + MEM[16290];
assign MEM[22060] = MEM[13416] + MEM[14656];
assign MEM[22061] = MEM[13417] + MEM[14447];
assign MEM[22062] = MEM[13421] + MEM[13602];
assign MEM[22063] = MEM[13423] + MEM[16530];
assign MEM[22064] = MEM[13424] + MEM[13506];
assign MEM[22065] = MEM[13424] + MEM[14927];
assign MEM[22066] = MEM[13425] + MEM[15701];
assign MEM[22067] = MEM[13428] + MEM[20240];
assign MEM[22068] = MEM[13435] + MEM[16124];
assign MEM[22069] = MEM[13449] + MEM[14200];
assign MEM[22070] = MEM[13449] + MEM[15432];
assign MEM[22071] = MEM[13450] + MEM[16386];
assign MEM[22072] = MEM[13451] + MEM[14163];
assign MEM[22073] = MEM[13452] + MEM[14415];
assign MEM[22074] = MEM[13455] + MEM[14223];
assign MEM[22075] = MEM[13471] + MEM[15003];
assign MEM[22076] = MEM[13473] + MEM[15687];
assign MEM[22077] = MEM[13479] + MEM[16672];
assign MEM[22078] = MEM[13483] + MEM[14365];
assign MEM[22079] = MEM[13487] + MEM[17832];
assign MEM[22080] = MEM[13488] + MEM[14704];
assign MEM[22081] = MEM[13493] + MEM[14395];
assign MEM[22082] = MEM[13495] + MEM[13582];
assign MEM[22083] = MEM[13495] + MEM[13642];
assign MEM[22084] = MEM[13496] + MEM[15050];
assign MEM[22085] = MEM[13497] + MEM[13906];
assign MEM[22086] = MEM[13498] + MEM[14298];
assign MEM[22087] = MEM[13500] + MEM[11367];
assign MEM[22088] = MEM[13502] + MEM[13514];
assign MEM[22089] = MEM[13506] + MEM[16721];
assign MEM[22090] = MEM[13508] + MEM[16106];
assign MEM[22091] = MEM[13510] + MEM[16149];
assign MEM[22092] = MEM[13512] + MEM[14778];
assign MEM[22093] = MEM[13513] + MEM[21371];
assign MEM[22094] = MEM[13514] + MEM[16382];
assign MEM[22095] = MEM[13515] + MEM[13851];
assign MEM[22096] = MEM[13522] + MEM[15879];
assign MEM[22097] = MEM[13523] + MEM[14064];
assign MEM[22098] = MEM[13533] + MEM[14470];
assign MEM[22099] = MEM[13536] + MEM[14017];
assign MEM[22100] = MEM[13539] + MEM[16380];
assign MEM[22101] = MEM[13542] + MEM[14777];
assign MEM[22102] = MEM[13543] + MEM[15880];
assign MEM[22103] = MEM[13546] + MEM[20422];
assign MEM[22104] = MEM[13553] + MEM[15858];
assign MEM[22105] = MEM[13556] + MEM[14374];
assign MEM[22106] = MEM[13572] + MEM[13988];
assign MEM[22107] = MEM[13573] + MEM[6954];
assign MEM[22108] = MEM[13581] + MEM[18825];
assign MEM[22109] = MEM[13587] + MEM[13599];
assign MEM[22110] = MEM[13589] + MEM[13809];
assign MEM[22111] = MEM[13605] + MEM[14976];
assign MEM[22112] = MEM[13608] + MEM[14105];
assign MEM[22113] = MEM[13608] + MEM[15949];
assign MEM[22114] = MEM[13609] + MEM[14122];
assign MEM[22115] = MEM[13612] + MEM[16139];
assign MEM[22116] = MEM[13614] + MEM[14445];
assign MEM[22117] = MEM[13617] + MEM[17036];
assign MEM[22118] = MEM[13620] + MEM[14227];
assign MEM[22119] = MEM[13623] + MEM[14851];
assign MEM[22120] = MEM[13624] + MEM[13881];
assign MEM[22121] = MEM[13624] + MEM[21296];
assign MEM[22122] = MEM[13625] + MEM[14532];
assign MEM[22123] = MEM[13633] + MEM[14199];
assign MEM[22124] = MEM[13634] + MEM[14043];
assign MEM[22125] = MEM[13636] + MEM[16123];
assign MEM[22126] = MEM[13640] + MEM[13889];
assign MEM[22127] = MEM[13642] + MEM[13722];
assign MEM[22128] = MEM[13649] + MEM[15251];
assign MEM[22129] = MEM[13651] + MEM[16344];
assign MEM[22130] = MEM[13653] + MEM[15934];
assign MEM[22131] = MEM[13657] + MEM[15117];
assign MEM[22132] = MEM[13658] + MEM[14700];
assign MEM[22133] = MEM[13659] + MEM[17421];
assign MEM[22134] = MEM[13662] + MEM[13883];
assign MEM[22135] = MEM[13662] + MEM[15419];
assign MEM[22136] = MEM[13665] + MEM[13678];
assign MEM[22137] = MEM[13665] + MEM[15198];
assign MEM[22138] = MEM[13668] + MEM[13822];
assign MEM[22139] = MEM[13677] + MEM[17145];
assign MEM[22140] = MEM[13680] + MEM[17162];
assign MEM[22141] = MEM[13681] + MEM[16218];
assign MEM[22142] = MEM[13683] + MEM[13807];
assign MEM[22143] = MEM[13685] + MEM[14479];
assign MEM[22144] = MEM[13687] + MEM[17076];
assign MEM[22145] = MEM[13694] + MEM[15195];
assign MEM[22146] = MEM[13697] + MEM[18231];
assign MEM[22147] = MEM[13701] + MEM[14206];
assign MEM[22148] = MEM[13701] + MEM[14801];
assign MEM[22149] = MEM[13703] + MEM[15143];
assign MEM[22150] = MEM[13711] + MEM[14027];
assign MEM[22151] = MEM[13713] + MEM[13977];
assign MEM[22152] = MEM[13719] + MEM[14208];
assign MEM[22153] = MEM[13719] + MEM[15262];
assign MEM[22154] = MEM[13724] + MEM[14021];
assign MEM[22155] = MEM[13729] + MEM[14033];
assign MEM[22156] = MEM[13739] + MEM[14202];
assign MEM[22157] = MEM[13739] + MEM[19412];
assign MEM[22158] = MEM[13745] + MEM[16677];
assign MEM[22159] = MEM[13746] + MEM[16219];
assign MEM[22160] = MEM[13747] + MEM[11930];
assign MEM[22161] = MEM[13751] + MEM[15253];
assign MEM[22162] = MEM[13753] + MEM[8372];
assign MEM[22163] = MEM[13755] + MEM[14537];
assign MEM[22164] = MEM[13757] + MEM[14138];
assign MEM[22165] = MEM[13758] + MEM[14659];
assign MEM[22166] = MEM[13759] + MEM[16803];
assign MEM[22167] = MEM[13765] + MEM[13989];
assign MEM[22168] = MEM[13772] + MEM[20559];
assign MEM[22169] = MEM[13775] + MEM[14311];
assign MEM[22170] = MEM[13776] + MEM[14275];
assign MEM[22171] = MEM[13776] + MEM[16710];
assign MEM[22172] = MEM[13781] + MEM[17015];
assign MEM[22173] = MEM[13793] + MEM[19030];
assign MEM[22174] = MEM[13794] + MEM[14233];
assign MEM[22175] = MEM[13797] + MEM[16570];
assign MEM[22176] = MEM[13800] + MEM[16278];
assign MEM[22177] = MEM[13803] + MEM[14066];
assign MEM[22178] = MEM[13805] + MEM[21260];
assign MEM[22179] = MEM[13806] + MEM[19739];
assign MEM[22180] = MEM[13808] + MEM[17600];
assign MEM[22181] = MEM[13816] + MEM[15989];
assign MEM[22182] = MEM[13821] + MEM[15314];
assign MEM[22183] = MEM[13830] + MEM[18966];
assign MEM[22184] = MEM[13831] + MEM[14502];
assign MEM[22185] = MEM[13832] + MEM[10150];
assign MEM[22186] = MEM[13838] + MEM[14735];
assign MEM[22187] = MEM[13840] + MEM[14906];
assign MEM[22188] = MEM[13841] + MEM[14290];
assign MEM[22189] = MEM[13848] + MEM[15821];
assign MEM[22190] = MEM[13852] + MEM[16586];
assign MEM[22191] = MEM[13853] + MEM[14035];
assign MEM[22192] = MEM[13855] + MEM[16748];
assign MEM[22193] = MEM[13859] + MEM[13877];
assign MEM[22194] = MEM[13862] + MEM[15075];
assign MEM[22195] = MEM[13865] + MEM[14077];
assign MEM[22196] = MEM[13869] + MEM[14299];
assign MEM[22197] = MEM[13871] + MEM[16082];
assign MEM[22198] = MEM[13872] + MEM[14134];
assign MEM[22199] = MEM[13873] + MEM[14252];
assign MEM[22200] = MEM[13876] + MEM[15158];
assign MEM[22201] = MEM[13884] + MEM[14366];
assign MEM[22202] = MEM[13885] + MEM[15205];
assign MEM[22203] = MEM[13888] + MEM[14396];
assign MEM[22204] = MEM[13892] + MEM[15438];
assign MEM[22205] = MEM[13894] + MEM[14934];
assign MEM[22206] = MEM[13896] + MEM[15658];
assign MEM[22207] = MEM[13898] + MEM[14995];
assign MEM[22208] = MEM[13907] + MEM[14368];
assign MEM[22209] = MEM[13910] + MEM[14722];
assign MEM[22210] = MEM[13914] + MEM[14518];
assign MEM[22211] = MEM[13917] + MEM[15145];
assign MEM[22212] = MEM[13922] + MEM[16232];
assign MEM[22213] = MEM[13924] + MEM[14552];
assign MEM[22214] = MEM[13925] + MEM[15194];
assign MEM[22215] = MEM[13928] + MEM[15105];
assign MEM[22216] = MEM[13929] + MEM[14256];
assign MEM[22217] = MEM[13933] + MEM[14379];
assign MEM[22218] = MEM[13934] + MEM[15699];
assign MEM[22219] = MEM[13937] + MEM[14554];
assign MEM[22220] = MEM[13940] + MEM[10049];
assign MEM[22221] = MEM[13941] + MEM[15371];
assign MEM[22222] = MEM[13942] + MEM[14770];
assign MEM[22223] = MEM[13944] + MEM[15401];
assign MEM[22224] = MEM[13951] + MEM[14520];
assign MEM[22225] = MEM[13953] + MEM[14699];
assign MEM[22226] = MEM[13956] + MEM[14222];
assign MEM[22227] = MEM[13957] + MEM[14356];
assign MEM[22228] = MEM[13960] + MEM[15247];
assign MEM[22229] = MEM[13961] + MEM[14022];
assign MEM[22230] = MEM[13965] + MEM[15781];
assign MEM[22231] = MEM[13966] + MEM[14286];
assign MEM[22232] = MEM[13967] + MEM[15681];
assign MEM[22233] = MEM[13971] + MEM[15170];
assign MEM[22234] = MEM[13974] + MEM[15346];
assign MEM[22235] = MEM[13975] + MEM[15076];
assign MEM[22236] = MEM[13978] + MEM[14515];
assign MEM[22237] = MEM[13981] + MEM[14407];
assign MEM[22238] = MEM[13984] + MEM[14053];
assign MEM[22239] = MEM[13987] + MEM[14070];
assign MEM[22240] = MEM[13991] + MEM[15147];
assign MEM[22241] = MEM[13995] + MEM[15175];
assign MEM[22242] = MEM[13997] + MEM[14127];
assign MEM[22243] = MEM[13998] + MEM[14969];
assign MEM[22244] = MEM[13999] + MEM[15475];
assign MEM[22245] = MEM[14000] + MEM[14220];
assign MEM[22246] = MEM[14001] + MEM[14684];
assign MEM[22247] = MEM[14002] + MEM[15082];
assign MEM[22248] = MEM[14003] + MEM[14455];
assign MEM[22249] = MEM[14004] + MEM[14442];
assign MEM[22250] = MEM[14005] + MEM[14563];
assign MEM[22251] = MEM[14010] + MEM[14082];
assign MEM[22252] = MEM[14011] + MEM[14393];
assign MEM[22253] = MEM[14014] + MEM[16714];
assign MEM[22254] = MEM[14018] + MEM[15732];
assign MEM[22255] = MEM[14028] + MEM[16127];
assign MEM[22256] = MEM[14029] + MEM[14098];
assign MEM[22257] = MEM[14037] + MEM[14067];
assign MEM[22258] = MEM[14038] + MEM[16129];
assign MEM[22259] = MEM[14039] + MEM[15162];
assign MEM[22260] = MEM[14042] + MEM[14478];
assign MEM[22261] = MEM[14044] + MEM[14313];
assign MEM[22262] = MEM[14058] + MEM[14614];
assign MEM[22263] = MEM[14059] + MEM[15042];
assign MEM[22264] = MEM[14062] + MEM[14523];
assign MEM[22265] = MEM[14068] + MEM[14885];
assign MEM[22266] = MEM[14071] + MEM[15579];
assign MEM[22267] = MEM[14075] + MEM[14960];
assign MEM[22268] = MEM[14076] + MEM[15293];
assign MEM[22269] = MEM[14083] + MEM[15324];
assign MEM[22270] = MEM[14089] + MEM[15009];
assign MEM[22271] = MEM[14090] + MEM[15470];
assign MEM[22272] = MEM[14091] + MEM[15259];
assign MEM[22273] = MEM[14092] + MEM[14701];
assign MEM[22274] = MEM[14093] + MEM[18183];
assign MEM[22275] = MEM[14096] + MEM[16404];
assign MEM[22276] = MEM[14102] + MEM[15573];
assign MEM[22277] = MEM[14107] + MEM[14754];
assign MEM[22278] = MEM[14111] + MEM[14946];
assign MEM[22279] = MEM[14112] + MEM[15309];
assign MEM[22280] = MEM[14118] + MEM[17450];
assign MEM[22281] = MEM[14124] + MEM[14129];
assign MEM[22282] = MEM[14126] + MEM[15040];
assign MEM[22283] = MEM[14132] + MEM[14270];
assign MEM[22284] = MEM[14135] + MEM[15448];
assign MEM[22285] = MEM[14136] + MEM[15282];
assign MEM[22286] = MEM[14137] + MEM[15029];
assign MEM[22287] = MEM[14141] + MEM[14631];
assign MEM[22288] = MEM[14143] + MEM[14260];
assign MEM[22289] = MEM[14145] + MEM[15906];
assign MEM[22290] = MEM[14146] + MEM[14856];
assign MEM[22291] = MEM[14152] + MEM[14490];
assign MEM[22292] = MEM[14153] + MEM[14473];
assign MEM[22293] = MEM[14159] + MEM[15337];
assign MEM[22294] = MEM[14160] + MEM[14284];
assign MEM[22295] = MEM[14167] + MEM[14792];
assign MEM[22296] = MEM[14169] + MEM[16201];
assign MEM[22297] = MEM[14170] + MEM[15255];
assign MEM[22298] = MEM[14177] + MEM[15335];
assign MEM[22299] = MEM[14179] + MEM[14835];
assign MEM[22300] = MEM[14180] + MEM[17359];
assign MEM[22301] = MEM[14181] + MEM[14386];
assign MEM[22302] = MEM[14185] + MEM[16505];
assign MEM[22303] = MEM[14189] + MEM[15363];
assign MEM[22304] = MEM[14190] + MEM[16220];
assign MEM[22305] = MEM[14194] + MEM[14655];
assign MEM[22306] = MEM[14212] + MEM[14485];
assign MEM[22307] = MEM[14213] + MEM[10243];
assign MEM[22308] = MEM[14225] + MEM[16716];
assign MEM[22309] = MEM[14234] + MEM[15883];
assign MEM[22310] = MEM[14236] + MEM[14582];
assign MEM[22311] = MEM[14240] + MEM[15450];
assign MEM[22312] = MEM[14241] + MEM[14634];
assign MEM[22313] = MEM[14249] + MEM[14881];
assign MEM[22314] = MEM[14257] + MEM[15597];
assign MEM[22315] = MEM[14280] + MEM[14397];
assign MEM[22316] = MEM[14289] + MEM[14330];
assign MEM[22317] = MEM[14292] + MEM[14566];
assign MEM[22318] = MEM[14293] + MEM[14897];
assign MEM[22319] = MEM[14302] + MEM[16155];
assign MEM[22320] = MEM[14305] + MEM[14426];
assign MEM[22321] = MEM[14314] + MEM[14820];
assign MEM[22322] = MEM[14316] + MEM[16398];
assign MEM[22323] = MEM[14317] + MEM[14816];
assign MEM[22324] = MEM[14318] + MEM[14862];
assign MEM[22325] = MEM[14319] + MEM[16199];
assign MEM[22326] = MEM[14321] + MEM[14605];
assign MEM[22327] = MEM[14322] + MEM[14665];
assign MEM[22328] = MEM[14323] + MEM[14411];
assign MEM[22329] = MEM[14325] + MEM[14392];
assign MEM[22330] = MEM[14326] + MEM[14623];
assign MEM[22331] = MEM[14328] + MEM[14729];
assign MEM[22332] = MEM[14333] + MEM[14487];
assign MEM[22333] = MEM[14334] + MEM[14456];
assign MEM[22334] = MEM[14337] + MEM[15225];
assign MEM[22335] = MEM[14340] + MEM[14717];
assign MEM[22336] = MEM[14342] + MEM[14643];
assign MEM[22337] = MEM[14343] + MEM[15806];
assign MEM[22338] = MEM[14346] + MEM[15035];
assign MEM[22339] = MEM[14347] + MEM[16312];
assign MEM[22340] = MEM[14354] + MEM[14653];
assign MEM[22341] = MEM[14358] + MEM[16859];
assign MEM[22342] = MEM[14359] + MEM[14632];
assign MEM[22343] = MEM[14361] + MEM[14584];
assign MEM[22344] = MEM[14363] + MEM[15585];
assign MEM[22345] = MEM[14370] + MEM[14610];
assign MEM[22346] = MEM[14371] + MEM[14687];
assign MEM[22347] = MEM[14373] + MEM[14568];
assign MEM[22348] = MEM[14378] + MEM[14925];
assign MEM[22349] = MEM[14381] + MEM[14535];
assign MEM[22350] = MEM[14394] + MEM[15629];
assign MEM[22351] = MEM[14400] + MEM[14494];
assign MEM[22352] = MEM[14401] + MEM[14430];
assign MEM[22353] = MEM[14405] + MEM[10377];
assign MEM[22354] = MEM[14409] + MEM[15604];
assign MEM[22355] = MEM[14410] + MEM[16351];
assign MEM[22356] = MEM[14419] + MEM[16184];
assign MEM[22357] = MEM[14421] + MEM[15397];
assign MEM[22358] = MEM[14422] + MEM[14697];
assign MEM[22359] = MEM[14423] + MEM[14843];
assign MEM[22360] = MEM[14425] + MEM[16873];
assign MEM[22361] = MEM[14428] + MEM[15362];
assign MEM[22362] = MEM[14437] + MEM[14580];
assign MEM[22363] = MEM[14440] + MEM[15063];
assign MEM[22364] = MEM[14441] + MEM[15283];
assign MEM[22365] = MEM[14443] + MEM[14932];
assign MEM[22366] = MEM[14446] + MEM[17865];
assign MEM[22367] = MEM[14460] + MEM[14874];
assign MEM[22368] = MEM[14461] + MEM[16120];
assign MEM[22369] = MEM[14463] + MEM[16089];
assign MEM[22370] = MEM[14467] + MEM[16093];
assign MEM[22371] = MEM[14469] + MEM[15240];
assign MEM[22372] = MEM[14471] + MEM[17255];
assign MEM[22373] = MEM[14475] + MEM[9837];
assign MEM[22374] = MEM[14477] + MEM[14489];
assign MEM[22375] = MEM[14483] + MEM[16318];
assign MEM[22376] = MEM[14484] + MEM[15295];
assign MEM[22377] = MEM[14491] + MEM[14500];
assign MEM[22378] = MEM[14493] + MEM[15976];
assign MEM[22379] = MEM[14499] + MEM[16877];
assign MEM[22380] = MEM[14508] + MEM[15467];
assign MEM[22381] = MEM[14509] + MEM[14578];
assign MEM[22382] = MEM[14510] + MEM[16511];
assign MEM[22383] = MEM[14511] + MEM[14649];
assign MEM[22384] = MEM[14521] + MEM[16360];
assign MEM[22385] = MEM[14525] + MEM[16227];
assign MEM[22386] = MEM[14526] + MEM[16669];
assign MEM[22387] = MEM[14527] + MEM[14819];
assign MEM[22388] = MEM[14529] + MEM[15737];
assign MEM[22389] = MEM[14534] + MEM[15224];
assign MEM[22390] = MEM[14536] + MEM[17236];
assign MEM[22391] = MEM[14538] + MEM[15084];
assign MEM[22392] = MEM[14539] + MEM[15632];
assign MEM[22393] = MEM[14540] + MEM[14847];
assign MEM[22394] = MEM[14543] + MEM[17224];
assign MEM[22395] = MEM[14545] + MEM[16256];
assign MEM[22396] = MEM[14546] + MEM[15411];
assign MEM[22397] = MEM[14550] + MEM[15376];
assign MEM[22398] = MEM[14555] + MEM[17377];
assign MEM[22399] = MEM[14557] + MEM[14888];
assign MEM[22400] = MEM[14558] + MEM[14972];
assign MEM[22401] = MEM[14560] + MEM[15051];
assign MEM[22402] = MEM[14562] + MEM[16037];
assign MEM[22403] = MEM[14569] + MEM[15341];
assign MEM[22404] = MEM[14570] + MEM[16002];
assign MEM[22405] = MEM[14579] + MEM[14677];
assign MEM[22406] = MEM[14581] + MEM[15791];
assign MEM[22407] = MEM[14583] + MEM[14876];
assign MEM[22408] = MEM[14586] + MEM[14909];
assign MEM[22409] = MEM[14591] + MEM[14931];
assign MEM[22410] = MEM[14592] + MEM[16172];
assign MEM[22411] = MEM[14593] + MEM[15526];
assign MEM[22412] = MEM[14601] + MEM[15758];
assign MEM[22413] = MEM[14602] + MEM[14818];
assign MEM[22414] = MEM[14603] + MEM[15124];
assign MEM[22415] = MEM[14604] + MEM[15643];
assign MEM[22416] = MEM[14606] + MEM[14730];
assign MEM[22417] = MEM[14609] + MEM[15131];
assign MEM[22418] = MEM[14611] + MEM[16308];
assign MEM[22419] = MEM[14615] + MEM[16974];
assign MEM[22420] = MEM[14616] + MEM[15101];
assign MEM[22421] = MEM[14618] + MEM[16083];
assign MEM[22422] = MEM[14620] + MEM[15279];
assign MEM[22423] = MEM[14627] + MEM[15312];
assign MEM[22424] = MEM[14637] + MEM[15339];
assign MEM[22425] = MEM[14639] + MEM[14652];
assign MEM[22426] = MEM[14650] + MEM[15345];
assign MEM[22427] = MEM[14658] + MEM[17142];
assign MEM[22428] = MEM[14664] + MEM[16295];
assign MEM[22429] = MEM[14666] + MEM[14911];
assign MEM[22430] = MEM[14671] + MEM[15261];
assign MEM[22431] = MEM[14676] + MEM[15028];
assign MEM[22432] = MEM[14680] + MEM[14737];
assign MEM[22433] = MEM[14682] + MEM[15365];
assign MEM[22434] = MEM[14689] + MEM[15981];
assign MEM[22435] = MEM[14690] + MEM[16822];
assign MEM[22436] = MEM[14692] + MEM[14783];
assign MEM[22437] = MEM[14693] + MEM[16016];
assign MEM[22438] = MEM[14695] + MEM[17343];
assign MEM[22439] = MEM[14706] + MEM[14947];
assign MEM[22440] = MEM[14707] + MEM[16343];
assign MEM[22441] = MEM[14710] + MEM[15690];
assign MEM[22442] = MEM[14711] + MEM[15088];
assign MEM[22443] = MEM[14714] + MEM[16827];
assign MEM[22444] = MEM[14715] + MEM[14721];
assign MEM[22445] = MEM[14718] + MEM[16136];
assign MEM[22446] = MEM[14719] + MEM[14720];
assign MEM[22447] = MEM[14727] + MEM[17414];
assign MEM[22448] = MEM[14732] + MEM[7193];
assign MEM[22449] = MEM[14733] + MEM[14834];
assign MEM[22450] = MEM[14734] + MEM[14767];
assign MEM[22451] = MEM[14738] + MEM[14823];
assign MEM[22452] = MEM[14739] + MEM[15289];
assign MEM[22453] = MEM[14741] + MEM[14786];
assign MEM[22454] = MEM[14743] + MEM[16292];
assign MEM[22455] = MEM[14749] + MEM[15179];
assign MEM[22456] = MEM[14757] + MEM[16038];
assign MEM[22457] = MEM[14760] + MEM[17695];
assign MEM[22458] = MEM[14761] + MEM[15109];
assign MEM[22459] = MEM[14762] + MEM[14973];
assign MEM[22460] = MEM[14765] + MEM[15197];
assign MEM[22461] = MEM[14769] + MEM[16578];
assign MEM[22462] = MEM[14773] + MEM[17666];
assign MEM[22463] = MEM[14775] + MEM[16749];
assign MEM[22464] = MEM[14785] + MEM[11415];
assign MEM[22465] = MEM[14788] + MEM[14838];
assign MEM[22466] = MEM[14791] + MEM[16222];
assign MEM[22467] = MEM[14794] + MEM[16357];
assign MEM[22468] = MEM[14795] + MEM[15323];
assign MEM[22469] = MEM[14797] + MEM[14844];
assign MEM[22470] = MEM[14802] + MEM[17120];
assign MEM[22471] = MEM[14803] + MEM[15011];
assign MEM[22472] = MEM[14806] + MEM[16041];
assign MEM[22473] = MEM[14808] + MEM[15551];
assign MEM[22474] = MEM[14814] + MEM[15462];
assign MEM[22475] = MEM[14817] + MEM[16072];
assign MEM[22476] = MEM[14825] + MEM[14959];
assign MEM[22477] = MEM[14826] + MEM[15241];
assign MEM[22478] = MEM[14831] + MEM[15216];
assign MEM[22479] = MEM[14832] + MEM[14877];
assign MEM[22480] = MEM[14837] + MEM[15464];
assign MEM[22481] = MEM[14841] + MEM[15306];
assign MEM[22482] = MEM[14842] + MEM[16300];
assign MEM[22483] = MEM[14846] + MEM[15550];
assign MEM[22484] = MEM[14850] + MEM[19382];
assign MEM[22485] = MEM[14863] + MEM[15654];
assign MEM[22486] = MEM[14864] + MEM[15529];
assign MEM[22487] = MEM[14865] + MEM[15574];
assign MEM[22488] = MEM[14866] + MEM[16903];
assign MEM[22489] = MEM[14869] + MEM[17117];
assign MEM[22490] = MEM[14875] + MEM[14237];
assign MEM[22491] = MEM[14878] + MEM[9882];
assign MEM[22492] = MEM[14879] + MEM[16161];
assign MEM[22493] = MEM[14884] + MEM[14929];
assign MEM[22494] = MEM[14887] + MEM[15347];
assign MEM[22495] = MEM[14892] + MEM[16430];
assign MEM[22496] = MEM[14894] + MEM[14907];
assign MEM[22497] = MEM[14904] + MEM[11206];
assign MEM[22498] = MEM[14915] + MEM[16637];
assign MEM[22499] = MEM[14916] + MEM[15652];
assign MEM[22500] = MEM[14917] + MEM[15662];
assign MEM[22501] = MEM[14919] + MEM[15469];
assign MEM[22502] = MEM[14926] + MEM[15825];
assign MEM[22503] = MEM[14933] + MEM[15044];
assign MEM[22504] = MEM[14935] + MEM[16208];
assign MEM[22505] = MEM[14937] + MEM[16942];
assign MEM[22506] = MEM[14938] + MEM[17100];
assign MEM[22507] = MEM[14940] + MEM[15039];
assign MEM[22508] = MEM[14950] + MEM[16428];
assign MEM[22509] = MEM[14953] + MEM[16269];
assign MEM[22510] = MEM[14954] + MEM[16328];
assign MEM[22511] = MEM[14957] + MEM[16230];
assign MEM[22512] = MEM[14964] + MEM[15267];
assign MEM[22513] = MEM[14965] + MEM[15850];
assign MEM[22514] = MEM[14971] + MEM[15177];
assign MEM[22515] = MEM[14974] + MEM[16108];
assign MEM[22516] = MEM[14978] + MEM[15125];
assign MEM[22517] = MEM[14981] + MEM[8485];
assign MEM[22518] = MEM[14984] + MEM[18786];
assign MEM[22519] = MEM[14988] + MEM[15290];
assign MEM[22520] = MEM[14989] + MEM[15838];
assign MEM[22521] = MEM[14994] + MEM[15960];
assign MEM[22522] = MEM[15001] + MEM[16030];
assign MEM[22523] = MEM[15007] + MEM[16014];
assign MEM[22524] = MEM[15008] + MEM[15421];
assign MEM[22525] = MEM[15013] + MEM[16488];
assign MEM[22526] = MEM[15018] + MEM[15169];
assign MEM[22527] = MEM[15038] + MEM[15118];
assign MEM[22528] = MEM[15048] + MEM[15121];
assign MEM[22529] = MEM[15052] + MEM[15260];
assign MEM[22530] = MEM[15053] + MEM[16024];
assign MEM[22531] = MEM[15054] + MEM[16980];
assign MEM[22532] = MEM[15058] + MEM[15387];
assign MEM[22533] = MEM[15059] + MEM[15146];
assign MEM[22534] = MEM[15064] + MEM[16905];
assign MEM[22535] = MEM[15068] + MEM[15349];
assign MEM[22536] = MEM[15069] + MEM[15528];
assign MEM[22537] = MEM[15074] + MEM[15275];
assign MEM[22538] = MEM[15078] + MEM[16297];
assign MEM[22539] = MEM[15079] + MEM[15353];
assign MEM[22540] = MEM[15086] + MEM[15454];
assign MEM[22541] = MEM[15090] + MEM[16032];
assign MEM[22542] = MEM[15095] + MEM[16946];
assign MEM[22543] = MEM[15097] + MEM[15343];
assign MEM[22544] = MEM[15107] + MEM[5203];
assign MEM[22545] = MEM[15113] + MEM[15457];
assign MEM[22546] = MEM[15119] + MEM[15779];
assign MEM[22547] = MEM[15120] + MEM[16352];
assign MEM[22548] = MEM[15132] + MEM[16182];
assign MEM[22549] = MEM[15135] + MEM[15413];
assign MEM[22550] = MEM[15138] + MEM[16574];
assign MEM[22551] = MEM[15139] + MEM[16503];
assign MEM[22552] = MEM[15142] + MEM[15212];
assign MEM[22553] = MEM[15153] + MEM[17301];
assign MEM[22554] = MEM[15155] + MEM[15824];
assign MEM[22555] = MEM[15164] + MEM[20933];
assign MEM[22556] = MEM[15173] + MEM[16678];
assign MEM[22557] = MEM[15174] + MEM[15917];
assign MEM[22558] = MEM[15181] + MEM[17886];
assign MEM[22559] = MEM[15186] + MEM[14905];
assign MEM[22560] = MEM[15187] + MEM[15229];
assign MEM[22561] = MEM[15188] + MEM[16639];
assign MEM[22562] = MEM[15189] + MEM[16132];
assign MEM[22563] = MEM[15199] + MEM[15898];
assign MEM[22564] = MEM[15206] + MEM[15956];
assign MEM[22565] = MEM[15207] + MEM[16732];
assign MEM[22566] = MEM[15208] + MEM[15593];
assign MEM[22567] = MEM[15213] + MEM[16323];
assign MEM[22568] = MEM[15222] + MEM[16941];
assign MEM[22569] = MEM[15223] + MEM[16243];
assign MEM[22570] = MEM[15231] + MEM[17137];
assign MEM[22571] = MEM[15233] + MEM[16998];
assign MEM[22572] = MEM[15234] + MEM[16885];
assign MEM[22573] = MEM[15239] + MEM[15263];
assign MEM[22574] = MEM[15246] + MEM[16122];
assign MEM[22575] = MEM[15252] + MEM[15287];
assign MEM[22576] = MEM[15258] + MEM[15610];
assign MEM[22577] = MEM[15265] + MEM[20345];
assign MEM[22578] = MEM[15273] + MEM[15683];
assign MEM[22579] = MEM[15276] + MEM[17215];
assign MEM[22580] = MEM[15278] + MEM[16519];
assign MEM[22581] = MEM[15284] + MEM[15486];
assign MEM[22582] = MEM[15294] + MEM[16248];
assign MEM[22583] = MEM[15297] + MEM[16730];
assign MEM[22584] = MEM[15299] + MEM[15015];
assign MEM[22585] = MEM[15302] + MEM[15418];
assign MEM[22586] = MEM[15303] + MEM[16241];
assign MEM[22587] = MEM[15305] + MEM[15518];
assign MEM[22588] = MEM[15308] + MEM[16498];
assign MEM[22589] = MEM[15311] + MEM[15490];
assign MEM[22590] = MEM[15315] + MEM[16613];
assign MEM[22591] = MEM[15322] + MEM[15919];
assign MEM[22592] = MEM[15328] + MEM[15773];
assign MEM[22593] = MEM[15329] + MEM[19089];
assign MEM[22594] = MEM[15331] + MEM[16869];
assign MEM[22595] = MEM[15338] + MEM[18483];
assign MEM[22596] = MEM[15348] + MEM[15549];
assign MEM[22597] = MEM[15354] + MEM[17747];
assign MEM[22598] = MEM[15355] + MEM[15941];
assign MEM[22599] = MEM[15366] + MEM[20222];
assign MEM[22600] = MEM[15369] + MEM[16728];
assign MEM[22601] = MEM[15373] + MEM[15430];
assign MEM[22602] = MEM[15375] + MEM[16359];
assign MEM[22603] = MEM[15378] + MEM[15947];
assign MEM[22604] = MEM[15384] + MEM[14807];
assign MEM[22605] = MEM[15389] + MEM[20890];
assign MEM[22606] = MEM[15392] + MEM[15530];
assign MEM[22607] = MEM[15395] + MEM[15697];
assign MEM[22608] = MEM[15396] + MEM[16494];
assign MEM[22609] = MEM[15399] + MEM[18049];
assign MEM[22610] = MEM[15402] + MEM[10015];
assign MEM[22611] = MEM[15406] + MEM[15456];
assign MEM[22612] = MEM[15410] + MEM[16464];
assign MEM[22613] = MEM[15415] + MEM[15416];
assign MEM[22614] = MEM[15422] + MEM[17164];
assign MEM[22615] = MEM[15423] + MEM[15849];
assign MEM[22616] = MEM[15429] + MEM[8105];
assign MEM[22617] = MEM[15433] + MEM[15613];
assign MEM[22618] = MEM[15437] + MEM[16372];
assign MEM[22619] = MEM[15439] + MEM[16447];
assign MEM[22620] = MEM[15442] + MEM[16459];
assign MEM[22621] = MEM[15443] + MEM[16281];
assign MEM[22622] = MEM[15444] + MEM[15481];
assign MEM[22623] = MEM[15449] + MEM[16109];
assign MEM[22624] = MEM[15451] + MEM[15768];
assign MEM[22625] = MEM[15463] + MEM[15943];
assign MEM[22626] = MEM[15468] + MEM[16440];
assign MEM[22627] = MEM[15474] + MEM[17426];
assign MEM[22628] = MEM[15478] + MEM[15644];
assign MEM[22629] = MEM[15479] + MEM[21210];
assign MEM[22630] = MEM[15483] + MEM[16515];
assign MEM[22631] = MEM[15487] + MEM[16886];
assign MEM[22632] = MEM[15492] + MEM[16433];
assign MEM[22633] = MEM[15494] + MEM[17039];
assign MEM[22634] = MEM[15496] + MEM[16554];
assign MEM[22635] = MEM[15497] + MEM[11201];
assign MEM[22636] = MEM[15500] + MEM[15575];
assign MEM[22637] = MEM[15517] + MEM[16062];
assign MEM[22638] = MEM[15524] + MEM[17165];
assign MEM[22639] = MEM[15537] + MEM[16235];
assign MEM[22640] = MEM[15538] + MEM[15586];
assign MEM[22641] = MEM[15553] + MEM[15969];
assign MEM[22642] = MEM[15557] + MEM[15885];
assign MEM[22643] = MEM[15559] + MEM[15998];
assign MEM[22644] = MEM[15560] + MEM[15722];
assign MEM[22645] = MEM[15561] + MEM[16437];
assign MEM[22646] = MEM[15569] + MEM[15686];
assign MEM[22647] = MEM[15577] + MEM[16830];
assign MEM[22648] = MEM[15589] + MEM[16480];
assign MEM[22649] = MEM[15594] + MEM[16153];
assign MEM[22650] = MEM[15603] + MEM[15671];
assign MEM[22651] = MEM[15611] + MEM[18367];
assign MEM[22652] = MEM[15618] + MEM[15763];
assign MEM[22653] = MEM[15620] + MEM[16681];
assign MEM[22654] = MEM[15622] + MEM[15747];
assign MEM[22655] = MEM[15626] + MEM[16898];
assign MEM[22656] = MEM[15653] + MEM[16050];
assign MEM[22657] = MEM[15668] + MEM[18438];
assign MEM[22658] = MEM[15693] + MEM[17131];
assign MEM[22659] = MEM[15696] + MEM[16019];
assign MEM[22660] = MEM[15703] + MEM[15864];
assign MEM[22661] = MEM[15705] + MEM[20831];
assign MEM[22662] = MEM[15709] + MEM[16125];
assign MEM[22663] = MEM[15712] + MEM[16467];
assign MEM[22664] = MEM[15714] + MEM[15435];
assign MEM[22665] = MEM[15718] + MEM[19059];
assign MEM[22666] = MEM[15719] + MEM[16186];
assign MEM[22667] = MEM[15727] + MEM[14451];
assign MEM[22668] = MEM[15736] + MEM[17393];
assign MEM[22669] = MEM[15741] + MEM[17191];
assign MEM[22670] = MEM[15751] + MEM[16641];
assign MEM[22671] = MEM[15754] + MEM[16154];
assign MEM[22672] = MEM[15765] + MEM[17256];
assign MEM[22673] = MEM[15766] + MEM[20274];
assign MEM[22674] = MEM[15767] + MEM[18885];
assign MEM[22675] = MEM[15777] + MEM[16416];
assign MEM[22676] = MEM[15792] + MEM[17366];
assign MEM[22677] = MEM[15812] + MEM[17242];
assign MEM[22678] = MEM[15828] + MEM[17108];
assign MEM[22679] = MEM[15829] + MEM[16687];
assign MEM[22680] = MEM[15832] + MEM[15996];
assign MEM[22681] = MEM[15837] + MEM[16522];
assign MEM[22682] = MEM[15839] + MEM[19639];
assign MEM[22683] = MEM[15846] + MEM[17182];
assign MEM[22684] = MEM[15854] + MEM[16745];
assign MEM[22685] = MEM[15863] + MEM[16141];
assign MEM[22686] = MEM[15866] + MEM[19201];
assign MEM[22687] = MEM[15869] + MEM[11647];
assign MEM[22688] = MEM[15873] + MEM[20046];
assign MEM[22689] = MEM[15874] + MEM[16679];
assign MEM[22690] = MEM[15878] + MEM[15913];
assign MEM[22691] = MEM[15887] + MEM[17710];
assign MEM[22692] = MEM[15889] + MEM[16616];
assign MEM[22693] = MEM[15890] + MEM[15144];
assign MEM[22694] = MEM[15894] + MEM[16391];
assign MEM[22695] = MEM[15904] + MEM[19482];
assign MEM[22696] = MEM[15912] + MEM[15122];
assign MEM[22697] = MEM[15922] + MEM[16789];
assign MEM[22698] = MEM[15926] + MEM[15851];
assign MEM[22699] = MEM[15954] + MEM[17757];
assign MEM[22700] = MEM[15955] + MEM[6478];
assign MEM[22701] = MEM[15959] + MEM[16395];
assign MEM[22702] = MEM[15961] + MEM[16406];
assign MEM[22703] = MEM[15973] + MEM[17004];
assign MEM[22704] = MEM[15978] + MEM[16329];
assign MEM[22705] = MEM[16006] + MEM[17384];
assign MEM[22706] = MEM[16010] + MEM[17030];
assign MEM[22707] = MEM[16011] + MEM[21618];
assign MEM[22708] = MEM[16012] + MEM[16107];
assign MEM[22709] = MEM[16022] + MEM[16077];
assign MEM[22710] = MEM[16029] + MEM[16370];
assign MEM[22711] = MEM[16043] + MEM[16336];
assign MEM[22712] = MEM[16045] + MEM[15580];
assign MEM[22713] = MEM[16048] + MEM[16673];
assign MEM[22714] = MEM[16056] + MEM[16205];
assign MEM[22715] = MEM[16067] + MEM[16378];
assign MEM[22716] = MEM[16075] + MEM[21806];
assign MEM[22717] = MEM[16098] + MEM[16920];
assign MEM[22718] = MEM[16099] + MEM[11577];
assign MEM[22719] = MEM[16100] + MEM[15209];
assign MEM[22720] = MEM[16101] + MEM[17348];
assign MEM[22721] = MEM[16114] + MEM[16251];
assign MEM[22722] = MEM[16115] + MEM[17208];
assign MEM[22723] = MEM[16133] + MEM[15485];
assign MEM[22724] = MEM[16135] + MEM[16507];
assign MEM[22725] = MEM[16146] + MEM[16709];
assign MEM[22726] = MEM[16159] + MEM[16763];
assign MEM[22727] = MEM[16173] + MEM[15564];
assign MEM[22728] = MEM[16179] + MEM[14993];
assign MEM[22729] = MEM[16202] + MEM[16712];
assign MEM[22730] = MEM[16204] + MEM[17453];
assign MEM[22731] = MEM[16229] + MEM[17371];
assign MEM[22732] = MEM[16237] + MEM[16888];
assign MEM[22733] = MEM[16238] + MEM[16684];
assign MEM[22734] = MEM[16264] + MEM[16853];
assign MEM[22735] = MEM[16270] + MEM[18007];
assign MEM[22736] = MEM[16288] + MEM[17287];
assign MEM[22737] = MEM[16299] + MEM[15706];
assign MEM[22738] = MEM[16305] + MEM[16482];
assign MEM[22739] = MEM[16306] + MEM[16979];
assign MEM[22740] = MEM[16315] + MEM[5333];
assign MEM[22741] = MEM[16319] + MEM[17098];
assign MEM[22742] = MEM[16325] + MEM[16583];
assign MEM[22743] = MEM[16337] + MEM[16593];
assign MEM[22744] = MEM[16353] + MEM[17295];
assign MEM[22745] = MEM[16365] + MEM[15842];
assign MEM[22746] = MEM[16374] + MEM[17309];
assign MEM[22747] = MEM[16383] + MEM[11413];
assign MEM[22748] = MEM[16396] + MEM[19693];
assign MEM[22749] = MEM[16405] + MEM[20880];
assign MEM[22750] = MEM[16407] + MEM[21581];
assign MEM[22751] = MEM[16408] + MEM[19823];
assign MEM[22752] = MEM[16421] + MEM[15522];
assign MEM[22753] = MEM[16431] + MEM[16461];
assign MEM[22754] = MEM[16435] + MEM[18664];
assign MEM[22755] = MEM[16443] + MEM[17077];
assign MEM[22756] = MEM[16444] + MEM[15628];
assign MEM[22757] = MEM[16449] + MEM[15608];
assign MEM[22758] = MEM[16451] + MEM[15480];
assign MEM[22759] = MEM[16453] + MEM[16854];
assign MEM[22760] = MEM[16455] + MEM[16706];
assign MEM[22761] = MEM[16457] + MEM[17011];
assign MEM[22762] = MEM[16463] + MEM[17157];
assign MEM[22763] = MEM[16477] + MEM[17240];
assign MEM[22764] = MEM[16485] + MEM[16615];
assign MEM[22765] = MEM[16486] + MEM[16322];
assign MEM[22766] = MEM[16490] + MEM[16871];
assign MEM[22767] = MEM[16495] + MEM[15990];
assign MEM[22768] = MEM[16497] + MEM[16567];
assign MEM[22769] = MEM[16543] + MEM[16524];
assign MEM[22770] = MEM[16564] + MEM[16909];
assign MEM[22771] = MEM[16572] + MEM[18824];
assign MEM[22772] = MEM[16580] + MEM[16910];
assign MEM[22773] = MEM[16582] + MEM[15350];
assign MEM[22774] = MEM[16590] + MEM[21219];
assign MEM[22775] = MEM[16596] + MEM[16356];
assign MEM[22776] = MEM[16597] + MEM[15708];
assign MEM[22777] = MEM[16608] + MEM[16110];
assign MEM[22778] = MEM[16609] + MEM[16758];
assign MEM[22779] = MEM[16610] + MEM[16629];
assign MEM[22780] = MEM[16623] + MEM[17210];
assign MEM[22781] = MEM[16633] + MEM[15698];
assign MEM[22782] = MEM[16635] + MEM[18956];
assign MEM[22783] = MEM[16647] + MEM[15081];
assign MEM[22784] = MEM[16659] + MEM[17303];
assign MEM[22785] = MEM[16661] + MEM[20245];
assign MEM[22786] = MEM[16671] + MEM[16977];
assign MEM[22787] = MEM[16688] + MEM[17629];
assign MEM[22788] = MEM[16697] + MEM[16489];
assign MEM[22789] = MEM[16713] + MEM[18715];
assign MEM[22790] = MEM[16722] + MEM[16837];
assign MEM[22791] = MEM[16744] + MEM[17213];
assign MEM[22792] = MEM[16751] + MEM[17174];
assign MEM[22793] = MEM[16753] + MEM[16213];
assign MEM[22794] = MEM[16761] + MEM[17168];
assign MEM[22795] = MEM[16765] + MEM[15843];
assign MEM[22796] = MEM[16770] + MEM[16646];
assign MEM[22797] = MEM[16772] + MEM[17001];
assign MEM[22798] = MEM[16775] + MEM[15546];
assign MEM[22799] = MEM[16782] + MEM[17623];
assign MEM[22800] = MEM[16797] + MEM[20168];
assign MEM[22801] = MEM[16801] + MEM[17119];
assign MEM[22802] = MEM[16805] + MEM[17448];
assign MEM[22803] = MEM[16806] + MEM[16214];
assign MEM[22804] = MEM[16811] + MEM[17044];
assign MEM[22805] = MEM[16820] + MEM[15584];
assign MEM[22806] = MEM[16824] + MEM[18166];
assign MEM[22807] = MEM[16841] + MEM[19878];
assign MEM[22808] = MEM[16845] + MEM[15488];
assign MEM[22809] = MEM[16851] + MEM[16313];
assign MEM[22810] = MEM[16861] + MEM[16604];
assign MEM[22811] = MEM[16862] + MEM[16039];
assign MEM[22812] = MEM[16882] + MEM[17193];
assign MEM[22813] = MEM[16883] + MEM[19140];
assign MEM[22814] = MEM[16889] + MEM[15383];
assign MEM[22815] = MEM[16890] + MEM[17178];
assign MEM[22816] = MEM[16893] + MEM[19916];
assign MEM[22817] = MEM[16895] + MEM[17645];
assign MEM[22818] = MEM[16897] + MEM[13905];
assign MEM[22819] = MEM[16900] + MEM[19395];
assign MEM[22820] = MEM[16901] + MEM[17151];
assign MEM[22821] = MEM[16924] + MEM[16415];
assign MEM[22822] = MEM[16925] + MEM[18936];
assign MEM[22823] = MEM[16928] + MEM[17229];
assign MEM[22824] = MEM[16933] + MEM[15980];
assign MEM[22825] = MEM[16934] + MEM[17249];
assign MEM[22826] = MEM[16937] + MEM[16410];
assign MEM[22827] = MEM[16944] + MEM[16843];
assign MEM[22828] = MEM[16950] + MEM[15805];
assign MEM[22829] = MEM[16960] + MEM[17025];
assign MEM[22830] = MEM[16964] + MEM[16198];
assign MEM[22831] = MEM[16970] + MEM[17270];
assign MEM[22832] = MEM[16971] + MEM[15720];
assign MEM[22833] = MEM[16981] + MEM[19271];
assign MEM[22834] = MEM[16991] + MEM[14184];
assign MEM[22835] = MEM[16995] + MEM[20271];
assign MEM[22836] = MEM[17005] + MEM[15986];
assign MEM[22837] = MEM[17018] + MEM[15971];
assign MEM[22838] = MEM[17027] + MEM[16000];
assign MEM[22839] = MEM[17031] + MEM[15595];
assign MEM[22840] = MEM[17034] + MEM[16558];
assign MEM[22841] = MEM[17037] + MEM[17163];
assign MEM[22842] = MEM[17040] + MEM[16649];
assign MEM[22843] = MEM[17043] + MEM[17839];
assign MEM[22844] = MEM[17059] + MEM[14731];
assign MEM[22845] = MEM[17064] + MEM[16719];
assign MEM[22846] = MEM[17069] + MEM[18629];
assign MEM[22847] = MEM[17071] + MEM[16148];
assign MEM[22848] = MEM[17078] + MEM[20785];
assign MEM[22849] = MEM[17094] + MEM[17258];
assign MEM[22850] = MEM[17103] + MEM[16429];
assign MEM[22851] = MEM[17106] + MEM[16071];
assign MEM[22852] = MEM[17109] + MEM[17386];
assign MEM[22853] = MEM[17110] + MEM[16849];
assign MEM[22854] = MEM[17111] + MEM[19108];
assign MEM[22855] = MEM[17112] + MEM[17340];
assign MEM[22856] = MEM[17140] + MEM[16725];
assign MEM[22857] = MEM[17159] + MEM[16948];
assign MEM[22858] = MEM[17172] + MEM[17375];
assign MEM[22859] = MEM[17194] + MEM[16327];
assign MEM[22860] = MEM[17196] + MEM[17336];
assign MEM[22861] = MEM[17199] + MEM[19950];
assign MEM[22862] = MEM[17225] + MEM[16747];
assign MEM[22863] = MEM[17230] + MEM[17976];
assign MEM[22864] = MEM[17234] + MEM[20460];
assign MEM[22865] = MEM[17235] + MEM[17374];
assign MEM[22866] = MEM[17248] + MEM[15540];
assign MEM[22867] = MEM[17252] + MEM[16800];
assign MEM[22868] = MEM[17253] + MEM[16619];
assign MEM[22869] = MEM[17261] + MEM[17866];
assign MEM[22870] = MEM[17291] + MEM[16951];
assign MEM[22871] = MEM[17300] + MEM[17662];
assign MEM[22872] = MEM[17306] + MEM[16802];
assign MEM[22873] = MEM[17317] + MEM[18773];
assign MEM[22874] = MEM[17321] + MEM[21436];
assign MEM[22875] = MEM[17331] + MEM[17160];
assign MEM[22876] = MEM[17342] + MEM[17074];
assign MEM[22877] = MEM[17344] + MEM[16371];
assign MEM[22878] = MEM[17347] + MEM[19623];
assign MEM[22879] = MEM[17350] + MEM[16674];
assign MEM[22880] = MEM[17360] + MEM[15679];
assign MEM[22881] = MEM[17372] + MEM[21348];
assign MEM[22882] = MEM[17389] + MEM[15508];
assign MEM[22883] = MEM[17390] + MEM[17732];
assign MEM[22884] = MEM[17413] + MEM[16993];
assign MEM[22885] = MEM[17415] + MEM[16528];
assign MEM[22886] = MEM[17433] + MEM[5670];
assign MEM[22887] = MEM[17464] + MEM[19226];
assign MEM[22888] = MEM[17471] + MEM[21127];
assign MEM[22889] = MEM[17472] + MEM[15682];
assign MEM[22890] = MEM[17482] + MEM[16984];
assign MEM[22891] = MEM[17485] + MEM[16581];
assign MEM[22892] = MEM[17488] + MEM[17048];
assign MEM[22893] = MEM[17529] + MEM[15185];
assign MEM[22894] = MEM[17534] + MEM[21103];
assign MEM[22895] = MEM[17535] + MEM[18902];
assign MEM[22896] = MEM[17539] + MEM[18816];
assign MEM[22897] = MEM[17559] + MEM[20749];
assign MEM[22898] = MEM[17563] + MEM[20923];
assign MEM[22899] = MEM[17565] + MEM[16556];
assign MEM[22900] = MEM[17567] + MEM[22033];
assign MEM[22901] = MEM[17573] + MEM[20649];
assign MEM[22902] = MEM[17585] + MEM[16675];
assign MEM[22903] = MEM[17602] + MEM[21324];
assign MEM[22904] = MEM[17625] + MEM[16119];
assign MEM[22905] = MEM[17627] + MEM[16134];
assign MEM[22906] = MEM[17667] + MEM[20857];
assign MEM[22907] = MEM[17693] + MEM[16303];
assign MEM[22908] = MEM[17696] + MEM[16793];
assign MEM[22909] = MEM[17709] + MEM[15588];
assign MEM[22910] = MEM[17716] + MEM[17226];
assign MEM[22911] = MEM[17723] + MEM[16887];
assign MEM[22912] = MEM[17740] + MEM[20681];
assign MEM[22913] = MEM[17742] + MEM[15161];
assign MEM[22914] = MEM[17754] + MEM[17469];
assign MEM[22915] = MEM[17756] + MEM[21430];
assign MEM[22916] = MEM[17758] + MEM[17381];
assign MEM[22917] = MEM[17759] + MEM[16260];
assign MEM[22918] = MEM[17769] + MEM[17293];
assign MEM[22919] = MEM[17782] + MEM[14297];
assign MEM[22920] = MEM[17786] + MEM[16017];
assign MEM[22921] = MEM[17796] + MEM[22013];
assign MEM[22922] = MEM[17799] + MEM[17973];
assign MEM[22923] = MEM[17806] + MEM[19835];
assign MEM[22924] = MEM[17813] + MEM[21871];
assign MEM[22925] = MEM[17822] + MEM[19425];
assign MEM[22926] = MEM[17827] + MEM[16676];
assign MEM[22927] = MEM[17850] + MEM[15830];
assign MEM[22928] = MEM[17861] + MEM[16347];
assign MEM[22929] = MEM[17864] + MEM[19585];
assign MEM[22930] = MEM[17868] + MEM[17148];
assign MEM[22931] = MEM[17877] + MEM[20954];
assign MEM[22932] = MEM[17884] + MEM[19010];
assign MEM[22933] = MEM[17888] + MEM[16321];
assign MEM[22934] = MEM[17894] + MEM[16537];
assign MEM[22935] = MEM[17902] + MEM[22258];
assign MEM[22936] = MEM[17903] + MEM[22293];
assign MEM[22937] = MEM[17905] + MEM[16051];
assign MEM[22938] = MEM[17907] + MEM[16054];
assign MEM[22939] = MEM[17911] + MEM[15739];
assign MEM[22940] = MEM[17921] + MEM[16663];
assign MEM[22941] = MEM[17923] + MEM[14188];
assign MEM[22942] = MEM[17930] + MEM[21598];
assign MEM[22943] = MEM[17935] + MEM[20863];
assign MEM[22944] = MEM[17937] + MEM[16216];
assign MEM[22945] = MEM[17977] + MEM[17367];
assign MEM[22946] = MEM[17979] + MEM[17023];
assign MEM[22947] = MEM[17992] + MEM[22564];
assign MEM[22948] = MEM[17996] + MEM[15493];
assign MEM[22949] = MEM[18004] + MEM[16599];
assign MEM[22950] = MEM[18017] + MEM[16664];
assign MEM[22951] = MEM[18020] + MEM[14766];
assign MEM[22952] = MEM[18028] + MEM[21895];
assign MEM[22953] = MEM[18069] + MEM[17026];
assign MEM[22954] = MEM[18079] + MEM[16417];
assign MEM[22955] = MEM[18081] + MEM[20714];
assign MEM[22956] = MEM[18082] + MEM[15523];
assign MEM[22957] = MEM[18089] + MEM[20561];
assign MEM[22958] = MEM[18108] + MEM[16496];
assign MEM[22959] = MEM[18109] + MEM[21394];
assign MEM[22960] = MEM[18120] + MEM[21841];
assign MEM[22961] = MEM[18124] + MEM[21453];
assign MEM[22962] = MEM[18132] + MEM[21790];
assign MEM[22963] = MEM[18139] + MEM[16812];
assign MEM[22964] = MEM[18143] + MEM[17335];
assign MEM[22965] = MEM[18147] + MEM[20363];
assign MEM[22966] = MEM[18148] + MEM[16349];
assign MEM[22967] = MEM[18151] + MEM[19956];
assign MEM[22968] = MEM[18155] + MEM[16655];
assign MEM[22969] = MEM[18158] + MEM[15721];
assign MEM[22970] = MEM[18195] + MEM[17177];
assign MEM[22971] = MEM[18210] + MEM[17265];
assign MEM[22972] = MEM[18223] + MEM[20294];
assign MEM[22973] = MEM[18240] + MEM[16508];
assign MEM[22974] = MEM[18243] + MEM[16209];
assign MEM[22975] = MEM[18254] + MEM[20921];
assign MEM[22976] = MEM[18255] + MEM[22295];
assign MEM[22977] = MEM[18258] + MEM[17316];
assign MEM[22978] = MEM[18261] + MEM[16298];
assign MEM[22979] = MEM[18265] + MEM[22300];
assign MEM[22980] = MEM[18307] + MEM[16832];
assign MEM[22981] = MEM[18315] + MEM[15884];
assign MEM[22982] = MEM[18316] + MEM[17275];
assign MEM[22983] = MEM[18319] + MEM[17288];
assign MEM[22984] = MEM[18325] + MEM[22084];
assign MEM[22985] = MEM[18333] + MEM[17022];
assign MEM[22986] = MEM[18340] + MEM[18363];
assign MEM[22987] = MEM[18344] + MEM[17459];
assign MEM[22988] = MEM[18352] + MEM[16930];
assign MEM[22989] = MEM[18358] + MEM[16682];
assign MEM[22990] = MEM[18361] + MEM[21026];
assign MEM[22991] = MEM[18372] + MEM[17396];
assign MEM[22992] = MEM[18388] + MEM[22511];
assign MEM[22993] = MEM[18389] + MEM[20673];
assign MEM[22994] = MEM[18413] + MEM[17216];
assign MEM[22995] = MEM[18429] + MEM[21955];
assign MEM[22996] = MEM[18436] + MEM[16475];
assign MEM[22997] = MEM[18441] + MEM[16852];
assign MEM[22998] = MEM[18444] + MEM[18941];
assign MEM[22999] = MEM[18447] + MEM[21164];
assign MEM[23000] = MEM[18453] + MEM[16693];
assign MEM[23001] = MEM[18454] + MEM[22746];
assign MEM[23002] = MEM[18457] + MEM[16804];
assign MEM[23003] = MEM[18462] + MEM[21645];
assign MEM[23004] = MEM[18474] + MEM[22407];
assign MEM[23005] = MEM[18476] + MEM[17289];
assign MEM[23006] = MEM[18498] + MEM[17167];
assign MEM[23007] = MEM[18500] + MEM[21070];
assign MEM[23008] = MEM[18503] + MEM[21801];
assign MEM[23009] = MEM[18507] + MEM[20059];
assign MEM[23010] = MEM[18517] + MEM[21762];
assign MEM[23011] = MEM[18521] + MEM[22652];
assign MEM[23012] = MEM[18526] + MEM[18863];
assign MEM[23013] = MEM[18539] + MEM[22725];
assign MEM[23014] = MEM[18558] + MEM[21607];
assign MEM[23015] = MEM[18559] + MEM[20433];
assign MEM[23016] = MEM[18583] + MEM[17232];
assign MEM[23017] = MEM[18590] + MEM[21418];
assign MEM[23018] = MEM[18591] + MEM[22600];
assign MEM[23019] = MEM[18593] + MEM[20547];
assign MEM[23020] = MEM[18598] + MEM[15554];
assign MEM[23021] = MEM[18599] + MEM[16975];
assign MEM[23022] = MEM[18607] + MEM[15870];
assign MEM[23023] = MEM[18609] + MEM[15809];
assign MEM[23024] = MEM[18610] + MEM[21958];
assign MEM[23025] = MEM[18616] + MEM[16735];
assign MEM[23026] = MEM[18617] + MEM[16042];
assign MEM[23027] = MEM[18623] + MEM[16896];
assign MEM[23028] = MEM[18636] + MEM[21381];
assign MEM[23029] = MEM[18646] + MEM[21856];
assign MEM[23030] = MEM[18672] + MEM[21449];
assign MEM[23031] = MEM[18674] + MEM[22417];
assign MEM[23032] = MEM[18689] + MEM[17281];
assign MEM[23033] = MEM[18696] + MEM[16792];
assign MEM[23034] = MEM[18700] + MEM[22655];
assign MEM[23035] = MEM[18708] + MEM[16829];
assign MEM[23036] = MEM[18718] + MEM[15966];
assign MEM[23037] = MEM[18738] + MEM[15619];
assign MEM[23038] = MEM[18758] + MEM[21457];
assign MEM[23039] = MEM[18762] + MEM[17397];
assign MEM[23040] = MEM[18772] + MEM[17408];
assign MEM[23041] = MEM[18790] + MEM[16899];
assign MEM[23042] = MEM[18799] + MEM[16988];
assign MEM[23043] = MEM[18800] + MEM[16445];
assign MEM[23044] = MEM[18810] + MEM[21570];
assign MEM[23045] = MEM[18815] + MEM[17314];
assign MEM[23046] = MEM[18839] + MEM[16717];
assign MEM[23047] = MEM[18846] + MEM[20696];
assign MEM[23048] = MEM[18849] + MEM[20784];
assign MEM[23049] = MEM[18855] + MEM[16990];
assign MEM[23050] = MEM[18891] + MEM[17130];
assign MEM[23051] = MEM[18895] + MEM[15738];
assign MEM[23052] = MEM[18899] + MEM[16947];
assign MEM[23053] = MEM[18903] + MEM[15304];
assign MEM[23054] = MEM[18905] + MEM[20598];
assign MEM[23055] = MEM[18911] + MEM[22849];
assign MEM[23056] = MEM[18921] + MEM[20770];
assign MEM[23057] = MEM[18926] + MEM[9078];
assign MEM[23058] = MEM[18927] + MEM[17128];
assign MEM[23059] = MEM[18942] + MEM[17186];
assign MEM[23060] = MEM[18948] + MEM[21558];
assign MEM[23061] = MEM[18958] + MEM[16720];
assign MEM[23062] = MEM[18970] + MEM[16922];
assign MEM[23063] = MEM[18972] + MEM[16557];
assign MEM[23064] = MEM[18975] + MEM[21305];
assign MEM[23065] = MEM[18985] + MEM[17271];
assign MEM[23066] = MEM[18987] + MEM[21354];
assign MEM[23067] = MEM[19005] + MEM[21331];
assign MEM[23068] = MEM[19034] + MEM[16332];
assign MEM[23069] = MEM[19040] + MEM[20021];
assign MEM[23070] = MEM[19045] + MEM[16923];
assign MEM[23071] = MEM[19051] + MEM[21294];
assign MEM[23072] = MEM[19061] + MEM[16969];
assign MEM[23073] = MEM[19075] + MEM[19895];
assign MEM[23074] = MEM[19081] + MEM[22736];
assign MEM[23075] = MEM[19082] + MEM[21640];
assign MEM[23076] = MEM[19091] + MEM[16152];
assign MEM[23077] = MEM[19098] + MEM[22000];
assign MEM[23078] = MEM[19116] + MEM[21867];
assign MEM[23079] = MEM[19130] + MEM[14625];
assign MEM[23080] = MEM[19143] + MEM[15460];
assign MEM[23081] = MEM[19150] + MEM[21229];
assign MEM[23082] = MEM[19152] + MEM[21970];
assign MEM[23083] = MEM[19155] + MEM[15370];
assign MEM[23084] = MEM[19171] + MEM[17324];
assign MEM[23085] = MEM[19178] + MEM[21304];
assign MEM[23086] = MEM[19183] + MEM[21774];
assign MEM[23087] = MEM[19211] + MEM[16413];
assign MEM[23088] = MEM[19225] + MEM[16387];
assign MEM[23089] = MEM[19228] + MEM[21766];
assign MEM[23090] = MEM[19236] + MEM[22003];
assign MEM[23091] = MEM[19239] + MEM[15817];
assign MEM[23092] = MEM[19242] + MEM[21989];
assign MEM[23093] = MEM[19244] + MEM[15614];
assign MEM[23094] = MEM[19250] + MEM[20414];
assign MEM[23095] = MEM[19263] + MEM[16858];
assign MEM[23096] = MEM[19275] + MEM[21484];
assign MEM[23097] = MEM[19276] + MEM[21939];
assign MEM[23098] = MEM[19296] + MEM[17079];
assign MEM[23099] = MEM[19319] + MEM[16291];
assign MEM[23100] = MEM[19320] + MEM[19357];
assign MEM[23101] = MEM[19336] + MEM[21376];
assign MEM[23102] = MEM[19341] + MEM[16348];
assign MEM[23103] = MEM[19342] + MEM[21894];
assign MEM[23104] = MEM[19343] + MEM[21906];
assign MEM[23105] = MEM[19355] + MEM[16626];
assign MEM[23106] = MEM[19359] + MEM[16589];
assign MEM[23107] = MEM[19371] + MEM[17062];
assign MEM[23108] = MEM[19403] + MEM[17357];
assign MEM[23109] = MEM[19409] + MEM[22762];
assign MEM[23110] = MEM[19414] + MEM[15318];
assign MEM[23111] = MEM[19415] + MEM[14923];
assign MEM[23112] = MEM[19437] + MEM[20259];
assign MEM[23113] = MEM[19439] + MEM[15918];
assign MEM[23114] = MEM[19441] + MEM[21110];
assign MEM[23115] = MEM[19445] + MEM[17394];
assign MEM[23116] = MEM[19463] + MEM[17073];
assign MEM[23117] = MEM[19478] + MEM[21862];
assign MEM[23118] = MEM[19479] + MEM[15583];
assign MEM[23119] = MEM[19483] + MEM[15797];
assign MEM[23120] = MEM[19497] + MEM[22357];
assign MEM[23121] = MEM[19535] + MEM[15605];
assign MEM[23122] = MEM[19545] + MEM[16931];
assign MEM[23123] = MEM[19558] + MEM[20772];
assign MEM[23124] = MEM[19564] + MEM[21055];
assign MEM[23125] = MEM[19566] + MEM[16689];
assign MEM[23126] = MEM[19573] + MEM[16180];
assign MEM[23127] = MEM[19575] + MEM[17454];
assign MEM[23128] = MEM[19588] + MEM[16591];
assign MEM[23129] = MEM[19596] + MEM[21724];
assign MEM[23130] = MEM[19600] + MEM[17468];
assign MEM[23131] = MEM[19604] + MEM[15651];
assign MEM[23132] = MEM[19628] + MEM[22703];
assign MEM[23133] = MEM[19637] + MEM[11344];
assign MEM[23134] = MEM[19638] + MEM[20752];
assign MEM[23135] = MEM[19642] + MEM[21363];
assign MEM[23136] = MEM[19672] + MEM[15642];
assign MEM[23137] = MEM[19677] + MEM[16053];
assign MEM[23138] = MEM[19689] + MEM[16913];
assign MEM[23139] = MEM[19690] + MEM[15556];
assign MEM[23140] = MEM[19700] + MEM[16379];
assign MEM[23141] = MEM[19705] + MEM[15862];
assign MEM[23142] = MEM[19706] + MEM[16254];
assign MEM[23143] = MEM[19743] + MEM[21825];
assign MEM[23144] = MEM[19764] + MEM[22680];
assign MEM[23145] = MEM[19787] + MEM[22761];
assign MEM[23146] = MEM[19789] + MEM[15600];
assign MEM[23147] = MEM[19796] + MEM[16144];
assign MEM[23148] = MEM[19799] + MEM[15726];
assign MEM[23149] = MEM[19801] + MEM[22345];
assign MEM[23150] = MEM[19811] + MEM[16271];
assign MEM[23151] = MEM[19821] + MEM[22341];
assign MEM[23152] = MEM[19828] + MEM[15783];
assign MEM[23153] = MEM[19832] + MEM[21687];
assign MEM[23154] = MEM[19837] + MEM[16756];
assign MEM[23155] = MEM[19838] + MEM[15511];
assign MEM[23156] = MEM[19843] + MEM[22181];
assign MEM[23157] = MEM[19846] + MEM[17107];
assign MEM[23158] = MEM[19848] + MEM[15933];
assign MEM[23159] = MEM[19856] + MEM[21236];
assign MEM[23160] = MEM[19865] + MEM[22288];
assign MEM[23161] = MEM[19880] + MEM[15958];
assign MEM[23162] = MEM[19886] + MEM[20176];
assign MEM[23163] = MEM[19900] + MEM[15250];
assign MEM[23164] = MEM[19902] + MEM[16692];
assign MEM[23165] = MEM[19915] + MEM[16375];
assign MEM[23166] = MEM[19948] + MEM[22627];
assign MEM[23167] = MEM[19961] + MEM[20775];
assign MEM[23168] = MEM[19972] + MEM[16079];
assign MEM[23169] = MEM[19998] + MEM[16972];
assign MEM[23170] = MEM[20029] + MEM[21108];
assign MEM[23171] = MEM[20033] + MEM[10346];
assign MEM[23172] = MEM[20035] + MEM[15710];
assign MEM[23173] = MEM[20056] + MEM[20455];
assign MEM[23174] = MEM[20057] + MEM[21242];
assign MEM[23175] = MEM[20061] + MEM[16724];
assign MEM[23176] = MEM[20066] + MEM[16622];
assign MEM[23177] = MEM[20069] + MEM[15694];
assign MEM[23178] = MEM[20085] + MEM[14728];
assign MEM[23179] = MEM[20090] + MEM[16625];
assign MEM[23180] = MEM[20118] + MEM[15256];
assign MEM[23181] = MEM[20122] + MEM[16245];
assign MEM[23182] = MEM[20130] + MEM[16261];
assign MEM[23183] = MEM[20131] + MEM[22730];
assign MEM[23184] = MEM[20147] + MEM[21924];
assign MEM[23185] = MEM[20186] + MEM[16373];
assign MEM[23186] = MEM[20189] + MEM[17380];
assign MEM[23187] = MEM[20202] + MEM[22442];
assign MEM[23188] = MEM[20204] + MEM[21307];
assign MEM[23189] = MEM[20215] + MEM[20373];
assign MEM[23190] = MEM[20218] + MEM[21463];
assign MEM[23191] = MEM[20221] + MEM[16231];
assign MEM[23192] = MEM[20225] + MEM[15545];
assign MEM[23193] = MEM[20236] + MEM[22425];
assign MEM[23194] = MEM[20242] + MEM[20494];
assign MEM[23195] = MEM[20244] + MEM[22713];
assign MEM[23196] = MEM[20247] + MEM[17247];
assign MEM[23197] = MEM[20265] + MEM[20716];
assign MEM[23198] = MEM[20280] + MEM[16757];
assign MEM[23199] = MEM[20297] + MEM[15730];
assign MEM[23200] = MEM[20304] + MEM[22118];
assign MEM[23201] = MEM[20314] + MEM[16550];
assign MEM[23202] = MEM[20325] + MEM[16696];
assign MEM[23203] = MEM[20349] + MEM[16090];
assign MEM[23204] = MEM[20351] + MEM[15818];
assign MEM[23205] = MEM[20376] + MEM[22633];
assign MEM[23206] = MEM[20421] + MEM[15881];
assign MEM[23207] = MEM[20428] + MEM[15997];
assign MEM[23208] = MEM[20441] + MEM[16130];
assign MEM[23209] = MEM[20446] + MEM[22702];
assign MEM[23210] = MEM[20473] + MEM[15957];
assign MEM[23211] = MEM[20478] + MEM[16618];
assign MEM[23212] = MEM[20481] + MEM[16479];
assign MEM[23213] = MEM[20491] + MEM[22419];
assign MEM[23214] = MEM[20495] + MEM[16617];
assign MEM[23215] = MEM[20508] + MEM[21886];
assign MEM[23216] = MEM[20516] + MEM[15641];
assign MEM[23217] = MEM[20521] + MEM[15794];
assign MEM[23218] = MEM[20535] + MEM[22772];
assign MEM[23219] = MEM[20536] + MEM[21136];
assign MEM[23220] = MEM[20550] + MEM[15740];
assign MEM[23221] = MEM[20557] + MEM[21934];
assign MEM[23222] = MEM[20558] + MEM[21195];
assign MEM[23223] = MEM[20575] + MEM[16193];
assign MEM[23224] = MEM[20584] + MEM[15905];
assign MEM[23225] = MEM[20609] + MEM[17141];
assign MEM[23226] = MEM[20622] + MEM[22883];
assign MEM[23227] = MEM[20640] + MEM[17217];
assign MEM[23228] = MEM[20657] + MEM[16828];
assign MEM[23229] = MEM[20664] + MEM[17189];
assign MEM[23230] = MEM[20671] + MEM[15970];
assign MEM[23231] = MEM[20682] + MEM[15744];
assign MEM[23232] = MEM[20693] + MEM[22665];
assign MEM[23233] = MEM[20694] + MEM[15536];
assign MEM[23234] = MEM[20699] + MEM[21787];
assign MEM[23235] = MEM[20706] + MEM[22562];
assign MEM[23236] = MEM[20737] + MEM[15695];
assign MEM[23237] = MEM[20742] + MEM[16304];
assign MEM[23238] = MEM[20761] + MEM[15616];
assign MEM[23239] = MEM[20764] + MEM[16835];
assign MEM[23240] = MEM[20765] + MEM[11452];
assign MEM[23241] = MEM[20768] + MEM[16881];
assign MEM[23242] = MEM[20780] + MEM[16523];
assign MEM[23243] = MEM[20782] + MEM[21765];
assign MEM[23244] = MEM[20786] + MEM[17274];
assign MEM[23245] = MEM[20795] + MEM[16834];
assign MEM[23246] = MEM[20812] + MEM[22580];
assign MEM[23247] = MEM[20815] + MEM[22509];
assign MEM[23248] = MEM[20817] + MEM[22438];
assign MEM[23249] = MEM[20845] + MEM[17144];
assign MEM[23250] = MEM[20847] + MEM[15896];
assign MEM[23251] = MEM[20858] + MEM[22019];
assign MEM[23252] = MEM[20860] + MEM[16506];
assign MEM[23253] = MEM[20893] + MEM[17066];
assign MEM[23254] = MEM[20916] + MEM[15855];
assign MEM[23255] = MEM[20955] + MEM[16983];
assign MEM[23256] = MEM[20965] + MEM[16121];
assign MEM[23257] = MEM[21007] + MEM[15815];
assign MEM[23258] = MEM[21027] + MEM[17000];
assign MEM[23259] = MEM[21037] + MEM[16874];
assign MEM[23260] = MEM[21058] + MEM[16346];
assign MEM[23261] = MEM[21061] + MEM[15928];
assign MEM[23262] = MEM[21066] + MEM[22741];
assign MEM[23263] = MEM[21067] + MEM[15892];
assign MEM[23264] = MEM[21076] + MEM[16982];
assign MEM[23265] = MEM[21091] + MEM[16118];
assign MEM[23266] = MEM[21095] + MEM[22692];
assign MEM[23267] = MEM[21096] + MEM[17047];
assign MEM[23268] = MEM[21100] + MEM[17241];
assign MEM[23269] = MEM[21104] + MEM[15836];
assign MEM[23270] = MEM[21107] + MEM[15977];
assign MEM[23271] = MEM[21181] + MEM[16191];
assign MEM[23272] = MEM[21227] + MEM[22651];
assign MEM[23273] = MEM[21248] + MEM[17070];
assign MEM[23274] = MEM[21255] + MEM[22446];
assign MEM[23275] = MEM[21264] + MEM[16512];
assign MEM[23276] = MEM[21295] + MEM[15532];
assign MEM[23277] = MEM[21303] + MEM[15782];
assign MEM[23278] = MEM[21311] + MEM[15833];
assign MEM[23279] = MEM[21313] + MEM[22510];
assign MEM[23280] = MEM[21322] + MEM[15472];
assign MEM[23281] = MEM[21329] + MEM[17341];
assign MEM[23282] = MEM[21341] + MEM[22368];
assign MEM[23283] = MEM[21353] + MEM[16080];
assign MEM[23284] = MEM[21372] + MEM[16005];
assign MEM[23285] = MEM[21386] + MEM[21909];
assign MEM[23286] = MEM[21404] + MEM[22869];
assign MEM[23287] = MEM[21428] + MEM[22569];
assign MEM[23288] = MEM[21445] + MEM[22229];
assign MEM[23289] = MEM[21465] + MEM[21627];
assign MEM[23290] = MEM[21473] + MEM[16653];
assign MEM[23291] = MEM[21504] + MEM[17345];
assign MEM[23292] = MEM[21517] + MEM[16658];
assign MEM[23293] = MEM[21530] + MEM[16310];
assign MEM[23294] = MEM[21536] + MEM[17277];
assign MEM[23295] = MEM[21538] + MEM[22196];
assign MEM[23296] = MEM[21547] + MEM[22670];
assign MEM[23297] = MEM[21571] + MEM[16594];
assign MEM[23298] = MEM[21590] + MEM[15678];
assign MEM[23299] = MEM[21595] + MEM[17259];
assign MEM[23300] = MEM[21596] + MEM[22661];
assign MEM[23301] = MEM[21633] + MEM[16545];
assign MEM[23302] = MEM[21642] + MEM[22313];
assign MEM[23303] = MEM[21647] + MEM[17127];
assign MEM[23304] = MEM[21683] + MEM[16063];
assign MEM[23305] = MEM[21713] + MEM[16341];
assign MEM[23306] = MEM[21718] + MEM[16466];
assign MEM[23307] = MEM[21722] + MEM[15755];
assign MEM[23308] = MEM[21731] + MEM[17219];
assign MEM[23309] = MEM[21732] + MEM[16727];
assign MEM[23310] = MEM[21755] + MEM[22238];
assign MEM[23311] = MEM[21798] + MEM[17089];
assign MEM[23312] = MEM[21802] + MEM[15623];
assign MEM[23313] = MEM[21832] + MEM[16462];
assign MEM[23314] = MEM[21920] + MEM[17175];
assign MEM[23315] = MEM[21925] + MEM[17223];
assign MEM[23316] = MEM[21927] + MEM[16707];
assign MEM[23317] = MEM[21971] + MEM[16774];
assign MEM[23318] = MEM[21977] + MEM[15972];
assign MEM[23319] = MEM[22008] + MEM[15280];
assign MEM[23320] = MEM[22012] + MEM[17400];
assign MEM[23321] = MEM[22016] + MEM[17410];
assign MEM[23322] = MEM[22023] + MEM[22514];
assign MEM[23323] = MEM[22034] + MEM[16715];
assign MEM[23324] = MEM[22097] + MEM[16131];
assign MEM[23325] = MEM[22110] + MEM[15902];
assign MEM[23326] = MEM[22112] + MEM[17455];
assign MEM[23327] = MEM[22119] + MEM[16236];
assign MEM[23328] = MEM[22131] + MEM[15822];
assign MEM[23329] = MEM[22142] + MEM[15982];
assign MEM[23330] = MEM[22148] + MEM[15525];
assign MEM[23331] = MEM[22149] + MEM[17156];
assign MEM[23332] = MEM[22150] + MEM[22553];
assign MEM[23333] = MEM[22170] + MEM[15796];
assign MEM[23334] = MEM[22184] + MEM[16844];
assign MEM[23335] = MEM[22199] + MEM[16592];
assign MEM[23336] = MEM[22203] + MEM[15789];
assign MEM[23337] = MEM[22227] + MEM[22576];
assign MEM[23338] = MEM[22231] + MEM[15811];
assign MEM[23339] = MEM[22264] + MEM[16529];
assign MEM[23340] = MEM[22268] + MEM[22835];
assign MEM[23341] = MEM[22283] + MEM[17049];
assign MEM[23342] = MEM[22317] + MEM[16880];
assign MEM[23343] = MEM[22327] + MEM[16705];
assign MEM[23344] = MEM[22349] + MEM[16385];
assign MEM[23345] = MEM[22369] + MEM[17320];
assign MEM[23346] = MEM[22374] + MEM[16680];
assign MEM[23347] = MEM[22398] + MEM[23243];
assign MEM[23348] = MEM[22420] + MEM[16074];
assign MEM[23349] = MEM[22449] + MEM[16491];
assign MEM[23350] = MEM[22468] + MEM[16092];
assign MEM[23351] = MEM[22475] + MEM[17444];
assign MEM[23352] = MEM[22515] + MEM[16726];
assign MEM[23353] = MEM[22552] + MEM[15659];
assign MEM[23354] = MEM[22575] + MEM[15509];
assign MEM[23355] = MEM[22586] + MEM[17188];
assign MEM[23356] = MEM[22617] + MEM[16553];
assign MEM[23357] = MEM[22623] + MEM[17362];
assign MEM[23358] = MEM[22625] + MEM[17302];
assign MEM[23359] = MEM[22642] + MEM[16333];
assign MEM[23360] = MEM[22709] + MEM[16468];
assign MEM[23361] = MEM[22710] + MEM[16472];
assign MEM[23362] = MEM[22721] + MEM[17105];
assign MEM[23363] = MEM[22766] + MEM[17138];
assign MEM[23364] = MEM[22784] + MEM[17351];
assign MEM[23365] = MEM[55] + MEM[794];
assign MEM[23366] = MEM[63] + MEM[13102];
assign MEM[23367] = MEM[85] + MEM[3805];
assign MEM[23368] = MEM[94] + MEM[759];
assign MEM[23369] = MEM[109] + MEM[10331];
assign MEM[23370] = MEM[110] + MEM[5959];
assign MEM[23371] = MEM[111] + MEM[2892];
assign MEM[23372] = MEM[118] + MEM[9941];
assign MEM[23373] = MEM[127] + MEM[5629];
assign MEM[23374] = MEM[142] + MEM[1016];
assign MEM[23375] = MEM[149] + MEM[5638];
assign MEM[23376] = MEM[151] + MEM[4043];
assign MEM[23377] = MEM[157] + MEM[7967];
assign MEM[23378] = MEM[159] + MEM[4394];
assign MEM[23379] = MEM[166] + MEM[2364];
assign MEM[23380] = MEM[173] + MEM[5306];
assign MEM[23381] = MEM[174] + MEM[4307];
assign MEM[23382] = MEM[207] + MEM[6774];
assign MEM[23383] = MEM[214] + MEM[1787];
assign MEM[23384] = MEM[221] + MEM[1350];
assign MEM[23385] = MEM[279] + MEM[14418];
assign MEM[23386] = MEM[299] + MEM[10971];
assign MEM[23387] = MEM[302] + MEM[8418];
assign MEM[23388] = MEM[307] + MEM[8541];
assign MEM[23389] = MEM[310] + MEM[4349];
assign MEM[23390] = MEM[314] + MEM[9310];
assign MEM[23391] = MEM[325] + MEM[6404];
assign MEM[23392] = MEM[326] + MEM[1871];
assign MEM[23393] = MEM[330] + MEM[11715];
assign MEM[23394] = MEM[340] + MEM[8390];
assign MEM[23395] = MEM[342] + MEM[1219];
assign MEM[23396] = MEM[379] + MEM[1725];
assign MEM[23397] = MEM[388] + MEM[1021];
assign MEM[23398] = MEM[389] + MEM[5196];
assign MEM[23399] = MEM[406] + MEM[1247];
assign MEM[23400] = MEM[421] + MEM[6481];
assign MEM[23401] = MEM[439] + MEM[10547];
assign MEM[23402] = MEM[445] + MEM[7391];
assign MEM[23403] = MEM[461] + MEM[1579];
assign MEM[23404] = MEM[469] + MEM[14641];
assign MEM[23405] = MEM[482] + MEM[5365];
assign MEM[23406] = MEM[485] + MEM[2375];
assign MEM[23407] = MEM[500] + MEM[1819];
assign MEM[23408] = MEM[501] + MEM[4167];
assign MEM[23409] = MEM[507] + MEM[3436];
assign MEM[23410] = MEM[515] + MEM[4971];
assign MEM[23411] = MEM[516] + MEM[4319];
assign MEM[23412] = MEM[522] + MEM[6947];
assign MEM[23413] = MEM[523] + MEM[2655];
assign MEM[23414] = MEM[524] + MEM[1207];
assign MEM[23415] = MEM[526] + MEM[13208];
assign MEM[23416] = MEM[533] + MEM[1189];
assign MEM[23417] = MEM[537] + MEM[4009];
assign MEM[23418] = MEM[542] + MEM[3127];
assign MEM[23419] = MEM[550] + MEM[11088];
assign MEM[23420] = MEM[554] + MEM[5199];
assign MEM[23421] = MEM[571] + MEM[3405];
assign MEM[23422] = MEM[575] + MEM[11749];
assign MEM[23423] = MEM[580] + MEM[643];
assign MEM[23424] = MEM[582] + MEM[4477];
assign MEM[23425] = MEM[584] + MEM[1628];
assign MEM[23426] = MEM[588] + MEM[5988];
assign MEM[23427] = MEM[591] + MEM[1018];
assign MEM[23428] = MEM[593] + MEM[948];
assign MEM[23429] = MEM[599] + MEM[981];
assign MEM[23430] = MEM[612] + MEM[9612];
assign MEM[23431] = MEM[614] + MEM[5582];
assign MEM[23432] = MEM[620] + MEM[5637];
assign MEM[23433] = MEM[622] + MEM[8330];
assign MEM[23434] = MEM[626] + MEM[2188];
assign MEM[23435] = MEM[638] + MEM[4155];
assign MEM[23436] = MEM[639] + MEM[1299];
assign MEM[23437] = MEM[639] + MEM[6445];
assign MEM[23438] = MEM[655] + MEM[1943];
assign MEM[23439] = MEM[663] + MEM[2885];
assign MEM[23440] = MEM[702] + MEM[2651];
assign MEM[23441] = MEM[716] + MEM[1039];
assign MEM[23442] = MEM[718] + MEM[6069];
assign MEM[23443] = MEM[726] + MEM[11345];
assign MEM[23444] = MEM[732] + MEM[6826];
assign MEM[23445] = MEM[735] + MEM[8797];
assign MEM[23446] = MEM[738] + MEM[11559];
assign MEM[23447] = MEM[742] + MEM[5503];
assign MEM[23448] = MEM[752] + MEM[7817];
assign MEM[23449] = MEM[754] + MEM[11071];
assign MEM[23450] = MEM[763] + MEM[1422];
assign MEM[23451] = MEM[764] + MEM[3725];
assign MEM[23452] = MEM[779] + MEM[6558];
assign MEM[23453] = MEM[780] + MEM[2506];
assign MEM[23454] = MEM[784] + MEM[9648];
assign MEM[23455] = MEM[786] + MEM[6433];
assign MEM[23456] = MEM[798] + MEM[13635];
assign MEM[23457] = MEM[811] + MEM[910];
assign MEM[23458] = MEM[818] + MEM[3509];
assign MEM[23459] = MEM[819] + MEM[2652];
assign MEM[23460] = MEM[831] + MEM[9023];
assign MEM[23461] = MEM[832] + MEM[12938];
assign MEM[23462] = MEM[835] + MEM[15408];
assign MEM[23463] = MEM[840] + MEM[2491];
assign MEM[23464] = MEM[852] + MEM[2718];
assign MEM[23465] = MEM[858] + MEM[5475];
assign MEM[23466] = MEM[859] + MEM[3230];
assign MEM[23467] = MEM[860] + MEM[8556];
assign MEM[23468] = MEM[867] + MEM[2323];
assign MEM[23469] = MEM[868] + MEM[3175];
assign MEM[23470] = MEM[871] + MEM[3629];
assign MEM[23471] = MEM[874] + MEM[1028];
assign MEM[23472] = MEM[876] + MEM[5222];
assign MEM[23473] = MEM[878] + MEM[7333];
assign MEM[23474] = MEM[879] + MEM[3442];
assign MEM[23475] = MEM[885] + MEM[8987];
assign MEM[23476] = MEM[895] + MEM[10252];
assign MEM[23477] = MEM[910] + MEM[5870];
assign MEM[23478] = MEM[916] + MEM[11901];
assign MEM[23479] = MEM[918] + MEM[3123];
assign MEM[23480] = MEM[926] + MEM[4166];
assign MEM[23481] = MEM[939] + MEM[1654];
assign MEM[23482] = MEM[942] + MEM[1365];
assign MEM[23483] = MEM[949] + MEM[10432];
assign MEM[23484] = MEM[955] + MEM[2628];
assign MEM[23485] = MEM[959] + MEM[5260];
assign MEM[23486] = MEM[965] + MEM[7861];
assign MEM[23487] = MEM[972] + MEM[10751];
assign MEM[23488] = MEM[973] + MEM[1469];
assign MEM[23489] = MEM[980] + MEM[7506];
assign MEM[23490] = MEM[995] + MEM[4850];
assign MEM[23491] = MEM[996] + MEM[1726];
assign MEM[23492] = MEM[998] + MEM[11087];
assign MEM[23493] = MEM[999] + MEM[5351];
assign MEM[23494] = MEM[1002] + MEM[6086];
assign MEM[23495] = MEM[1003] + MEM[1371];
assign MEM[23496] = MEM[1005] + MEM[3555];
assign MEM[23497] = MEM[1007] + MEM[13387];
assign MEM[23498] = MEM[1018] + MEM[6294];
assign MEM[23499] = MEM[1026] + MEM[6682];
assign MEM[23500] = MEM[1029] + MEM[1451];
assign MEM[23501] = MEM[1035] + MEM[8566];
assign MEM[23502] = MEM[1036] + MEM[1182];
assign MEM[23503] = MEM[1047] + MEM[8399];
assign MEM[23504] = MEM[1054] + MEM[1851];
assign MEM[23505] = MEM[1059] + MEM[11840];
assign MEM[23506] = MEM[1079] + MEM[1302];
assign MEM[23507] = MEM[1127] + MEM[3743];
assign MEM[23508] = MEM[1157] + MEM[2102];
assign MEM[23509] = MEM[1157] + MEM[10129];
assign MEM[23510] = MEM[1162] + MEM[7275];
assign MEM[23511] = MEM[1166] + MEM[1754];
assign MEM[23512] = MEM[1173] + MEM[4355];
assign MEM[23513] = MEM[1175] + MEM[6023];
assign MEM[23514] = MEM[1191] + MEM[4411];
assign MEM[23515] = MEM[1196] + MEM[6538];
assign MEM[23516] = MEM[1203] + MEM[8461];
assign MEM[23517] = MEM[1211] + MEM[4965];
assign MEM[23518] = MEM[1212] + MEM[12734];
assign MEM[23519] = MEM[1213] + MEM[10178];
assign MEM[23520] = MEM[1220] + MEM[2029];
assign MEM[23521] = MEM[1230] + MEM[1327];
assign MEM[23522] = MEM[1234] + MEM[1452];
assign MEM[23523] = MEM[1236] + MEM[4325];
assign MEM[23524] = MEM[1244] + MEM[3374];
assign MEM[23525] = MEM[1254] + MEM[5813];
assign MEM[23526] = MEM[1258] + MEM[7072];
assign MEM[23527] = MEM[1274] + MEM[9902];
assign MEM[23528] = MEM[1275] + MEM[9933];
assign MEM[23529] = MEM[1276] + MEM[8266];
assign MEM[23530] = MEM[1282] + MEM[9913];
assign MEM[23531] = MEM[1284] + MEM[2402];
assign MEM[23532] = MEM[1310] + MEM[12857];
assign MEM[23533] = MEM[1314] + MEM[8757];
assign MEM[23534] = MEM[1317] + MEM[12040];
assign MEM[23535] = MEM[1326] + MEM[10237];
assign MEM[23536] = MEM[1341] + MEM[2084];
assign MEM[23537] = MEM[1364] + MEM[1890];
assign MEM[23538] = MEM[1366] + MEM[2103];
assign MEM[23539] = MEM[1373] + MEM[8446];
assign MEM[23540] = MEM[1378] + MEM[2804];
assign MEM[23541] = MEM[1382] + MEM[4295];
assign MEM[23542] = MEM[1383] + MEM[10567];
assign MEM[23543] = MEM[1389] + MEM[13206];
assign MEM[23544] = MEM[1395] + MEM[4739];
assign MEM[23545] = MEM[1397] + MEM[3359];
assign MEM[23546] = MEM[1407] + MEM[3022];
assign MEM[23547] = MEM[1415] + MEM[7218];
assign MEM[23548] = MEM[1430] + MEM[2499];
assign MEM[23549] = MEM[1438] + MEM[10862];
assign MEM[23550] = MEM[1443] + MEM[6323];
assign MEM[23551] = MEM[1447] + MEM[3443];
assign MEM[23552] = MEM[1451] + MEM[13920];
assign MEM[23553] = MEM[1463] + MEM[4565];
assign MEM[23554] = MEM[1474] + MEM[7356];
assign MEM[23555] = MEM[1476] + MEM[9447];
assign MEM[23556] = MEM[1483] + MEM[10868];
assign MEM[23557] = MEM[1486] + MEM[6708];
assign MEM[23558] = MEM[1492] + MEM[11566];
assign MEM[23559] = MEM[1494] + MEM[11629];
assign MEM[23560] = MEM[1499] + MEM[1935];
assign MEM[23561] = MEM[1500] + MEM[5010];
assign MEM[23562] = MEM[1509] + MEM[2996];
assign MEM[23563] = MEM[1515] + MEM[10541];
assign MEM[23564] = MEM[1518] + MEM[5250];
assign MEM[23565] = MEM[1525] + MEM[8349];
assign MEM[23566] = MEM[1548] + MEM[7336];
assign MEM[23567] = MEM[1550] + MEM[3221];
assign MEM[23568] = MEM[1567] + MEM[3614];
assign MEM[23569] = MEM[1575] + MEM[8033];
assign MEM[23570] = MEM[1597] + MEM[4087];
assign MEM[23571] = MEM[1604] + MEM[10594];
assign MEM[23572] = MEM[1643] + MEM[10359];
assign MEM[23573] = MEM[1669] + MEM[2566];
assign MEM[23574] = MEM[1670] + MEM[1750];
assign MEM[23575] = MEM[1674] + MEM[8899];
assign MEM[23576] = MEM[1675] + MEM[6651];
assign MEM[23577] = MEM[1677] + MEM[3403];
assign MEM[23578] = MEM[1708] + MEM[11879];
assign MEM[23579] = MEM[1716] + MEM[3236];
assign MEM[23580] = MEM[1722] + MEM[8191];
assign MEM[23581] = MEM[1741] + MEM[8648];
assign MEM[23582] = MEM[1744] + MEM[3003];
assign MEM[23583] = MEM[1749] + MEM[4381];
assign MEM[23584] = MEM[1755] + MEM[2612];
assign MEM[23585] = MEM[1770] + MEM[2326];
assign MEM[23586] = MEM[1772] + MEM[7249];
assign MEM[23587] = MEM[1778] + MEM[2279];
assign MEM[23588] = MEM[1788] + MEM[12476];
assign MEM[23589] = MEM[1797] + MEM[2171];
assign MEM[23590] = MEM[1798] + MEM[3967];
assign MEM[23591] = MEM[1799] + MEM[4292];
assign MEM[23592] = MEM[1806] + MEM[8000];
assign MEM[23593] = MEM[1810] + MEM[2971];
assign MEM[23594] = MEM[1831] + MEM[3469];
assign MEM[23595] = MEM[1845] + MEM[5748];
assign MEM[23596] = MEM[1854] + MEM[11221];
assign MEM[23597] = MEM[1855] + MEM[6302];
assign MEM[23598] = MEM[1862] + MEM[5671];
assign MEM[23599] = MEM[1876] + MEM[11807];
assign MEM[23600] = MEM[1892] + MEM[9396];
assign MEM[23601] = MEM[1893] + MEM[2141];
assign MEM[23602] = MEM[1894] + MEM[10942];
assign MEM[23603] = MEM[1898] + MEM[6143];
assign MEM[23604] = MEM[1900] + MEM[7087];
assign MEM[23605] = MEM[1901] + MEM[7977];
assign MEM[23606] = MEM[1908] + MEM[9906];
assign MEM[23607] = MEM[1918] + MEM[12860];
assign MEM[23608] = MEM[1923] + MEM[5094];
assign MEM[23609] = MEM[1930] + MEM[11017];
assign MEM[23610] = MEM[1934] + MEM[2827];
assign MEM[23611] = MEM[1942] + MEM[4092];
assign MEM[23612] = MEM[1949] + MEM[7520];
assign MEM[23613] = MEM[1955] + MEM[6724];
assign MEM[23614] = MEM[1999] + MEM[2960];
assign MEM[23615] = MEM[2003] + MEM[3047];
assign MEM[23616] = MEM[2005] + MEM[5183];
assign MEM[23617] = MEM[2006] + MEM[3314];
assign MEM[23618] = MEM[2007] + MEM[12661];
assign MEM[23619] = MEM[2020] + MEM[2907];
assign MEM[23620] = MEM[2021] + MEM[8192];
assign MEM[23621] = MEM[2038] + MEM[5550];
assign MEM[23622] = MEM[2051] + MEM[14337];
assign MEM[23623] = MEM[2058] + MEM[10027];
assign MEM[23624] = MEM[2068] + MEM[5762];
assign MEM[23625] = MEM[2071] + MEM[4551];
assign MEM[23626] = MEM[2074] + MEM[10068];
assign MEM[23627] = MEM[2094] + MEM[2631];
assign MEM[23628] = MEM[2106] + MEM[7708];
assign MEM[23629] = MEM[2107] + MEM[7518];
assign MEM[23630] = MEM[2111] + MEM[7762];
assign MEM[23631] = MEM[2114] + MEM[2556];
assign MEM[23632] = MEM[2115] + MEM[10451];
assign MEM[23633] = MEM[2117] + MEM[7528];
assign MEM[23634] = MEM[2118] + MEM[2378];
assign MEM[23635] = MEM[2123] + MEM[10389];
assign MEM[23636] = MEM[2127] + MEM[3431];
assign MEM[23637] = MEM[2133] + MEM[9743];
assign MEM[23638] = MEM[2134] + MEM[6901];
assign MEM[23639] = MEM[2136] + MEM[3279];
assign MEM[23640] = MEM[2142] + MEM[4683];
assign MEM[23641] = MEM[2149] + MEM[3620];
assign MEM[23642] = MEM[2162] + MEM[2470];
assign MEM[23643] = MEM[2180] + MEM[2444];
assign MEM[23644] = MEM[2181] + MEM[8469];
assign MEM[23645] = MEM[2182] + MEM[7877];
assign MEM[23646] = MEM[2190] + MEM[13281];
assign MEM[23647] = MEM[2206] + MEM[5717];
assign MEM[23648] = MEM[2208] + MEM[6739];
assign MEM[23649] = MEM[2213] + MEM[4189];
assign MEM[23650] = MEM[2214] + MEM[6812];
assign MEM[23651] = MEM[2217] + MEM[14602];
assign MEM[23652] = MEM[2220] + MEM[10477];
assign MEM[23653] = MEM[2223] + MEM[8223];
assign MEM[23654] = MEM[2229] + MEM[11443];
assign MEM[23655] = MEM[2236] + MEM[3237];
assign MEM[23656] = MEM[2251] + MEM[9505];
assign MEM[23657] = MEM[2258] + MEM[8881];
assign MEM[23658] = MEM[2263] + MEM[8617];
assign MEM[23659] = MEM[2268] + MEM[12144];
assign MEM[23660] = MEM[2269] + MEM[4858];
assign MEM[23661] = MEM[2277] + MEM[6194];
assign MEM[23662] = MEM[2291] + MEM[12088];
assign MEM[23663] = MEM[2295] + MEM[4158];
assign MEM[23664] = MEM[2301] + MEM[4695];
assign MEM[23665] = MEM[2302] + MEM[3664];
assign MEM[23666] = MEM[2303] + MEM[5900];
assign MEM[23667] = MEM[2307] + MEM[9661];
assign MEM[23668] = MEM[2308] + MEM[3716];
assign MEM[23669] = MEM[2311] + MEM[3797];
assign MEM[23670] = MEM[2312] + MEM[4729];
assign MEM[23671] = MEM[2325] + MEM[6854];
assign MEM[23672] = MEM[2341] + MEM[10917];
assign MEM[23673] = MEM[2346] + MEM[10600];
assign MEM[23674] = MEM[2357] + MEM[7771];
assign MEM[23675] = MEM[2359] + MEM[4826];
assign MEM[23676] = MEM[2360] + MEM[3213];
assign MEM[23677] = MEM[2370] + MEM[7878];
assign MEM[23678] = MEM[2391] + MEM[4883];
assign MEM[23679] = MEM[2398] + MEM[6955];
assign MEM[23680] = MEM[2404] + MEM[4669];
assign MEM[23681] = MEM[2410] + MEM[11423];
assign MEM[23682] = MEM[2416] + MEM[3853];
assign MEM[23683] = MEM[2421] + MEM[6583];
assign MEM[23684] = MEM[2428] + MEM[10964];
assign MEM[23685] = MEM[2430] + MEM[11265];
assign MEM[23686] = MEM[2432] + MEM[6213];
assign MEM[23687] = MEM[2435] + MEM[7374];
assign MEM[23688] = MEM[2441] + MEM[10168];
assign MEM[23689] = MEM[2443] + MEM[4475];
assign MEM[23690] = MEM[2453] + MEM[8146];
assign MEM[23691] = MEM[2454] + MEM[10113];
assign MEM[23692] = MEM[2459] + MEM[3391];
assign MEM[23693] = MEM[2483] + MEM[9668];
assign MEM[23694] = MEM[2494] + MEM[8871];
assign MEM[23695] = MEM[2495] + MEM[10647];
assign MEM[23696] = MEM[2498] + MEM[10424];
assign MEM[23697] = MEM[2516] + MEM[8007];
assign MEM[23698] = MEM[2519] + MEM[10182];
assign MEM[23699] = MEM[2523] + MEM[8276];
assign MEM[23700] = MEM[2534] + MEM[3628];
assign MEM[23701] = MEM[2542] + MEM[8501];
assign MEM[23702] = MEM[2546] + MEM[10315];
assign MEM[23703] = MEM[2547] + MEM[6132];
assign MEM[23704] = MEM[2548] + MEM[6062];
assign MEM[23705] = MEM[2549] + MEM[6142];
assign MEM[23706] = MEM[2550] + MEM[12053];
assign MEM[23707] = MEM[2551] + MEM[7393];
assign MEM[23708] = MEM[2557] + MEM[2726];
assign MEM[23709] = MEM[2563] + MEM[5991];
assign MEM[23710] = MEM[2578] + MEM[11963];
assign MEM[23711] = MEM[2581] + MEM[8753];
assign MEM[23712] = MEM[2582] + MEM[7167];
assign MEM[23713] = MEM[2583] + MEM[5043];
assign MEM[23714] = MEM[2587] + MEM[5356];
assign MEM[23715] = MEM[2596] + MEM[3835];
assign MEM[23716] = MEM[2619] + MEM[3166];
assign MEM[23717] = MEM[2635] + MEM[7738];
assign MEM[23718] = MEM[2636] + MEM[4522];
assign MEM[23719] = MEM[2639] + MEM[10890];
assign MEM[23720] = MEM[2643] + MEM[9661];
assign MEM[23721] = MEM[2644] + MEM[3707];
assign MEM[23722] = MEM[2648] + MEM[5676];
assign MEM[23723] = MEM[2656] + MEM[9256];
assign MEM[23724] = MEM[2657] + MEM[3035];
assign MEM[23725] = MEM[2658] + MEM[14767];
assign MEM[23726] = MEM[2660] + MEM[8715];
assign MEM[23727] = MEM[2662] + MEM[9691];
assign MEM[23728] = MEM[2666] + MEM[3421];
assign MEM[23729] = MEM[2667] + MEM[5839];
assign MEM[23730] = MEM[2670] + MEM[12676];
assign MEM[23731] = MEM[2674] + MEM[8769];
assign MEM[23732] = MEM[2675] + MEM[9624];
assign MEM[23733] = MEM[2678] + MEM[8249];
assign MEM[23734] = MEM[2686] + MEM[6133];
assign MEM[23735] = MEM[2695] + MEM[3668];
assign MEM[23736] = MEM[2711] + MEM[8055];
assign MEM[23737] = MEM[2720] + MEM[3821];
assign MEM[23738] = MEM[2722] + MEM[11627];
assign MEM[23739] = MEM[2723] + MEM[9213];
assign MEM[23740] = MEM[2738] + MEM[3052];
assign MEM[23741] = MEM[2739] + MEM[6417];
assign MEM[23742] = MEM[2747] + MEM[2948];
assign MEM[23743] = MEM[2748] + MEM[8387];
assign MEM[23744] = MEM[2749] + MEM[10685];
assign MEM[23745] = MEM[2752] + MEM[4468];
assign MEM[23746] = MEM[2763] + MEM[7271];
assign MEM[23747] = MEM[2767] + MEM[4630];
assign MEM[23748] = MEM[2770] + MEM[10937];
assign MEM[23749] = MEM[2771] + MEM[7450];
assign MEM[23750] = MEM[2772] + MEM[9647];
assign MEM[23751] = MEM[2776] + MEM[2968];
assign MEM[23752] = MEM[2778] + MEM[5316];
assign MEM[23753] = MEM[2798] + MEM[5434];
assign MEM[23754] = MEM[2812] + MEM[3717];
assign MEM[23755] = MEM[2815] + MEM[3396];
assign MEM[23756] = MEM[2819] + MEM[4691];
assign MEM[23757] = MEM[2831] + MEM[11772];
assign MEM[23758] = MEM[2835] + MEM[10894];
assign MEM[23759] = MEM[2869] + MEM[11524];
assign MEM[23760] = MEM[2870] + MEM[10056];
assign MEM[23761] = MEM[2932] + MEM[3922];
assign MEM[23762] = MEM[2939] + MEM[9112];
assign MEM[23763] = MEM[2955] + MEM[3234];
assign MEM[23764] = MEM[2957] + MEM[12735];
assign MEM[23765] = MEM[2962] + MEM[6707];
assign MEM[23766] = MEM[2963] + MEM[3895];
assign MEM[23767] = MEM[2973] + MEM[10982];
assign MEM[23768] = MEM[2974] + MEM[4179];
assign MEM[23769] = MEM[2976] + MEM[3242];
assign MEM[23770] = MEM[2981] + MEM[5519];
assign MEM[23771] = MEM[2987] + MEM[7005];
assign MEM[23772] = MEM[2989] + MEM[4060];
assign MEM[23773] = MEM[2997] + MEM[3590];
assign MEM[23774] = MEM[3014] + MEM[9584];
assign MEM[23775] = MEM[3020] + MEM[10739];
assign MEM[23776] = MEM[3023] + MEM[9072];
assign MEM[23777] = MEM[3046] + MEM[4718];
assign MEM[23778] = MEM[3053] + MEM[10255];
assign MEM[23779] = MEM[3061] + MEM[8998];
assign MEM[23780] = MEM[3063] + MEM[9717];
assign MEM[23781] = MEM[3084] + MEM[5053];
assign MEM[23782] = MEM[3090] + MEM[3562];
assign MEM[23783] = MEM[3091] + MEM[5070];
assign MEM[23784] = MEM[3102] + MEM[8620];
assign MEM[23785] = MEM[3110] + MEM[4235];
assign MEM[23786] = MEM[3118] + MEM[4143];
assign MEM[23787] = MEM[3124] + MEM[9462];
assign MEM[23788] = MEM[3126] + MEM[11831];
assign MEM[23789] = MEM[3143] + MEM[12444];
assign MEM[23790] = MEM[3174] + MEM[9684];
assign MEM[23791] = MEM[3189] + MEM[17620];
assign MEM[23792] = MEM[3195] + MEM[6804];
assign MEM[23793] = MEM[3200] + MEM[10923];
assign MEM[23794] = MEM[3218] + MEM[4293];
assign MEM[23795] = MEM[3219] + MEM[10492];
assign MEM[23796] = MEM[3226] + MEM[8782];
assign MEM[23797] = MEM[3229] + MEM[10733];
assign MEM[23798] = MEM[3235] + MEM[10396];
assign MEM[23799] = MEM[3238] + MEM[6297];
assign MEM[23800] = MEM[3243] + MEM[10434];
assign MEM[23801] = MEM[3254] + MEM[10021];
assign MEM[23802] = MEM[3261] + MEM[8381];
assign MEM[23803] = MEM[3283] + MEM[4126];
assign MEM[23804] = MEM[3284] + MEM[6486];
assign MEM[23805] = MEM[3290] + MEM[7334];
assign MEM[23806] = MEM[3292] + MEM[6489];
assign MEM[23807] = MEM[3295] + MEM[7911];
assign MEM[23808] = MEM[3300] + MEM[7117];
assign MEM[23809] = MEM[3306] + MEM[3486];
assign MEM[23810] = MEM[3334] + MEM[4946];
assign MEM[23811] = MEM[3341] + MEM[8756];
assign MEM[23812] = MEM[3366] + MEM[7093];
assign MEM[23813] = MEM[3367] + MEM[5983];
assign MEM[23814] = MEM[3407] + MEM[10279];
assign MEM[23815] = MEM[3412] + MEM[10856];
assign MEM[23816] = MEM[3413] + MEM[4726];
assign MEM[23817] = MEM[3428] + MEM[3623];
assign MEM[23818] = MEM[3434] + MEM[12667];
assign MEM[23819] = MEM[3445] + MEM[8434];
assign MEM[23820] = MEM[3450] + MEM[5764];
assign MEM[23821] = MEM[3454] + MEM[6864];
assign MEM[23822] = MEM[3463] + MEM[3476];
assign MEM[23823] = MEM[3474] + MEM[15067];
assign MEM[23824] = MEM[3485] + MEM[6363];
assign MEM[23825] = MEM[3498] + MEM[7147];
assign MEM[23826] = MEM[3508] + MEM[7689];
assign MEM[23827] = MEM[3510] + MEM[3605];
assign MEM[23828] = MEM[3522] + MEM[5069];
assign MEM[23829] = MEM[3530] + MEM[18094];
assign MEM[23830] = MEM[3538] + MEM[6644];
assign MEM[23831] = MEM[3551] + MEM[6669];
assign MEM[23832] = MEM[3558] + MEM[8135];
assign MEM[23833] = MEM[3574] + MEM[7695];
assign MEM[23834] = MEM[3579] + MEM[10855];
assign MEM[23835] = MEM[3599] + MEM[5942];
assign MEM[23836] = MEM[3611] + MEM[4997];
assign MEM[23837] = MEM[3626] + MEM[7596];
assign MEM[23838] = MEM[3632] + MEM[3640];
assign MEM[23839] = MEM[3636] + MEM[13721];
assign MEM[23840] = MEM[3643] + MEM[7790];
assign MEM[23841] = MEM[3648] + MEM[3904];
assign MEM[23842] = MEM[3652] + MEM[5591];
assign MEM[23843] = MEM[3655] + MEM[5668];
assign MEM[23844] = MEM[3656] + MEM[12231];
assign MEM[23845] = MEM[3661] + MEM[8340];
assign MEM[23846] = MEM[3666] + MEM[6117];
assign MEM[23847] = MEM[3672] + MEM[6635];
assign MEM[23848] = MEM[3674] + MEM[5037];
assign MEM[23849] = MEM[3691] + MEM[6021];
assign MEM[23850] = MEM[3694] + MEM[10452];
assign MEM[23851] = MEM[3730] + MEM[5402];
assign MEM[23852] = MEM[3733] + MEM[4989];
assign MEM[23853] = MEM[3735] + MEM[9064];
assign MEM[23854] = MEM[3743] + MEM[11251];
assign MEM[23855] = MEM[3747] + MEM[16394];
assign MEM[23856] = MEM[3750] + MEM[5389];
assign MEM[23857] = MEM[3755] + MEM[5382];
assign MEM[23858] = MEM[3763] + MEM[10721];
assign MEM[23859] = MEM[3764] + MEM[12828];
assign MEM[23860] = MEM[3773] + MEM[12102];
assign MEM[23861] = MEM[3782] + MEM[5548];
assign MEM[23862] = MEM[3786] + MEM[6322];
assign MEM[23863] = MEM[3794] + MEM[13330];
assign MEM[23864] = MEM[3795] + MEM[5953];
assign MEM[23865] = MEM[3799] + MEM[4750];
assign MEM[23866] = MEM[3806] + MEM[4471];
assign MEM[23867] = MEM[3822] + MEM[4429];
assign MEM[23868] = MEM[3826] + MEM[9909];
assign MEM[23869] = MEM[3831] + MEM[11534];
assign MEM[23870] = MEM[3834] + MEM[4851];
assign MEM[23871] = MEM[3842] + MEM[10271];
assign MEM[23872] = MEM[3847] + MEM[4909];
assign MEM[23873] = MEM[3852] + MEM[7549];
assign MEM[23874] = MEM[3861] + MEM[10529];
assign MEM[23875] = MEM[3871] + MEM[3901];
assign MEM[23876] = MEM[3876] + MEM[5541];
assign MEM[23877] = MEM[3877] + MEM[12121];
assign MEM[23878] = MEM[3880] + MEM[7135];
assign MEM[23879] = MEM[3882] + MEM[5770];
assign MEM[23880] = MEM[3883] + MEM[10292];
assign MEM[23881] = MEM[3884] + MEM[5313];
assign MEM[23882] = MEM[3900] + MEM[6246];
assign MEM[23883] = MEM[3902] + MEM[4287];
assign MEM[23884] = MEM[3918] + MEM[5556];
assign MEM[23885] = MEM[3924] + MEM[10146];
assign MEM[23886] = MEM[3931] + MEM[7098];
assign MEM[23887] = MEM[3933] + MEM[4410];
assign MEM[23888] = MEM[3940] + MEM[12993];
assign MEM[23889] = MEM[3943] + MEM[12356];
assign MEM[23890] = MEM[3947] + MEM[8947];
assign MEM[23891] = MEM[3949] + MEM[7723];
assign MEM[23892] = MEM[3957] + MEM[11034];
assign MEM[23893] = MEM[3962] + MEM[7460];
assign MEM[23894] = MEM[3965] + MEM[7411];
assign MEM[23895] = MEM[3974] + MEM[6746];
assign MEM[23896] = MEM[3987] + MEM[12321];
assign MEM[23897] = MEM[3994] + MEM[5653];
assign MEM[23898] = MEM[4003] + MEM[4050];
assign MEM[23899] = MEM[4020] + MEM[5013];
assign MEM[23900] = MEM[4046] + MEM[5915];
assign MEM[23901] = MEM[4047] + MEM[8120];
assign MEM[23902] = MEM[4059] + MEM[16538];
assign MEM[23903] = MEM[4062] + MEM[12108];
assign MEM[23904] = MEM[4078] + MEM[10611];
assign MEM[23905] = MEM[4091] + MEM[11583];
assign MEM[23906] = MEM[4098] + MEM[9454];
assign MEM[23907] = MEM[4101] + MEM[6348];
assign MEM[23908] = MEM[4103] + MEM[9970];
assign MEM[23909] = MEM[4107] + MEM[6928];
assign MEM[23910] = MEM[4111] + MEM[8874];
assign MEM[23911] = MEM[4128] + MEM[12757];
assign MEM[23912] = MEM[4132] + MEM[5727];
assign MEM[23913] = MEM[4141] + MEM[8973];
assign MEM[23914] = MEM[4146] + MEM[10508];
assign MEM[23915] = MEM[4151] + MEM[6367];
assign MEM[23916] = MEM[4156] + MEM[9097];
assign MEM[23917] = MEM[4162] + MEM[8742];
assign MEM[23918] = MEM[4163] + MEM[10786];
assign MEM[23919] = MEM[4165] + MEM[11273];
assign MEM[23920] = MEM[4172] + MEM[11805];
assign MEM[23921] = MEM[4187] + MEM[7881];
assign MEM[23922] = MEM[4189] + MEM[6740];
assign MEM[23923] = MEM[4206] + MEM[7800];
assign MEM[23924] = MEM[4214] + MEM[4229];
assign MEM[23925] = MEM[4228] + MEM[8219];
assign MEM[23926] = MEM[4246] + MEM[6389];
assign MEM[23927] = MEM[4251] + MEM[4285];
assign MEM[23928] = MEM[4252] + MEM[5268];
assign MEM[23929] = MEM[4262] + MEM[6949];
assign MEM[23930] = MEM[4271] + MEM[7331];
assign MEM[23931] = MEM[4291] + MEM[6749];
assign MEM[23932] = MEM[4292] + MEM[6562];
assign MEM[23933] = MEM[4300] + MEM[7660];
assign MEM[23934] = MEM[4309] + MEM[11570];
assign MEM[23935] = MEM[4310] + MEM[10802];
assign MEM[23936] = MEM[4315] + MEM[11926];
assign MEM[23937] = MEM[4316] + MEM[6649];
assign MEM[23938] = MEM[4318] + MEM[4511];
assign MEM[23939] = MEM[4324] + MEM[8385];
assign MEM[23940] = MEM[4335] + MEM[11321];
assign MEM[23941] = MEM[4350] + MEM[8502];
assign MEM[23942] = MEM[4359] + MEM[4439];
assign MEM[23943] = MEM[4359] + MEM[9853];
assign MEM[23944] = MEM[4363] + MEM[5230];
assign MEM[23945] = MEM[4372] + MEM[9712];
assign MEM[23946] = MEM[4380] + MEM[5772];
assign MEM[23947] = MEM[4399] + MEM[6729];
assign MEM[23948] = MEM[4402] + MEM[13236];
assign MEM[23949] = MEM[4405] + MEM[4770];
assign MEM[23950] = MEM[4407] + MEM[5005];
assign MEM[23951] = MEM[4412] + MEM[9631];
assign MEM[23952] = MEM[4418] + MEM[6404];
assign MEM[23953] = MEM[4420] + MEM[8653];
assign MEM[23954] = MEM[4427] + MEM[5188];
assign MEM[23955] = MEM[4435] + MEM[5206];
assign MEM[23956] = MEM[4442] + MEM[13547];
assign MEM[23957] = MEM[4447] + MEM[9658];
assign MEM[23958] = MEM[4460] + MEM[6312];
assign MEM[23959] = MEM[4461] + MEM[4927];
assign MEM[23960] = MEM[4466] + MEM[11924];
assign MEM[23961] = MEM[4469] + MEM[7325];
assign MEM[23962] = MEM[4479] + MEM[11456];
assign MEM[23963] = MEM[4486] + MEM[4722];
assign MEM[23964] = MEM[4487] + MEM[4557];
assign MEM[23965] = MEM[4493] + MEM[5542];
assign MEM[23966] = MEM[4508] + MEM[10202];
assign MEM[23967] = MEM[4509] + MEM[7977];
assign MEM[23968] = MEM[4517] + MEM[10268];
assign MEM[23969] = MEM[4525] + MEM[12541];
assign MEM[23970] = MEM[4531] + MEM[6637];
assign MEM[23971] = MEM[4542] + MEM[7548];
assign MEM[23972] = MEM[4548] + MEM[10052];
assign MEM[23973] = MEM[4558] + MEM[4967];
assign MEM[23974] = MEM[4562] + MEM[4796];
assign MEM[23975] = MEM[4564] + MEM[14556];
assign MEM[23976] = MEM[4567] + MEM[5903];
assign MEM[23977] = MEM[4573] + MEM[8558];
assign MEM[23978] = MEM[4582] + MEM[7763];
assign MEM[23979] = MEM[4583] + MEM[11899];
assign MEM[23980] = MEM[4587] + MEM[8217];
assign MEM[23981] = MEM[4595] + MEM[7718];
assign MEM[23982] = MEM[4605] + MEM[13641];
assign MEM[23983] = MEM[4623] + MEM[10718];
assign MEM[23984] = MEM[4635] + MEM[10210];
assign MEM[23985] = MEM[4651] + MEM[5917];
assign MEM[23986] = MEM[4658] + MEM[6354];
assign MEM[23987] = MEM[4659] + MEM[11938];
assign MEM[23988] = MEM[4676] + MEM[5815];
assign MEM[23989] = MEM[4693] + MEM[9359];
assign MEM[23990] = MEM[4715] + MEM[7128];
assign MEM[23991] = MEM[4742] + MEM[16065];
assign MEM[23992] = MEM[4743] + MEM[9871];
assign MEM[23993] = MEM[4767] + MEM[7442];
assign MEM[23994] = MEM[4772] + MEM[6038];
assign MEM[23995] = MEM[4780] + MEM[5771];
assign MEM[23996] = MEM[4782] + MEM[11910];
assign MEM[23997] = MEM[4805] + MEM[12688];
assign MEM[23998] = MEM[4813] + MEM[14374];
assign MEM[23999] = MEM[4819] + MEM[6664];
assign MEM[24000] = MEM[4820] + MEM[10018];
assign MEM[24001] = MEM[4838] + MEM[8279];
assign MEM[24002] = MEM[4842] + MEM[9674];
assign MEM[24003] = MEM[4852] + MEM[11587];
assign MEM[24004] = MEM[4855] + MEM[12817];
assign MEM[24005] = MEM[4867] + MEM[6306];
assign MEM[24006] = MEM[4868] + MEM[12116];
assign MEM[24007] = MEM[4869] + MEM[7389];
assign MEM[24008] = MEM[4871] + MEM[5678];
assign MEM[24009] = MEM[4876] + MEM[9277];
assign MEM[24010] = MEM[4887] + MEM[4916];
assign MEM[24011] = MEM[4911] + MEM[6270];
assign MEM[24012] = MEM[4915] + MEM[6568];
assign MEM[24013] = MEM[4917] + MEM[9034];
assign MEM[24014] = MEM[4949] + MEM[5253];
assign MEM[24015] = MEM[4950] + MEM[13998];
assign MEM[24016] = MEM[4962] + MEM[7324];
assign MEM[24017] = MEM[4966] + MEM[9398];
assign MEM[24018] = MEM[4972] + MEM[14848];
assign MEM[24019] = MEM[4973] + MEM[10421];
assign MEM[24020] = MEM[4987] + MEM[7863];
assign MEM[24021] = MEM[5003] + MEM[5471];
assign MEM[24022] = MEM[5006] + MEM[8361];
assign MEM[24023] = MEM[5007] + MEM[6380];
assign MEM[24024] = MEM[5019] + MEM[6172];
assign MEM[24025] = MEM[5021] + MEM[12874];
assign MEM[24026] = MEM[5023] + MEM[5098];
assign MEM[24027] = MEM[5026] + MEM[8822];
assign MEM[24028] = MEM[5031] + MEM[12695];
assign MEM[24029] = MEM[5038] + MEM[10895];
assign MEM[24030] = MEM[5046] + MEM[11562];
assign MEM[24031] = MEM[5068] + MEM[8775];
assign MEM[24032] = MEM[5075] + MEM[6204];
assign MEM[24033] = MEM[5083] + MEM[8019];
assign MEM[24034] = MEM[5084] + MEM[7533];
assign MEM[24035] = MEM[5087] + MEM[6933];
assign MEM[24036] = MEM[5091] + MEM[6946];
assign MEM[24037] = MEM[5094] + MEM[11863];
assign MEM[24038] = MEM[5111] + MEM[9531];
assign MEM[24039] = MEM[5115] + MEM[7286];
assign MEM[24040] = MEM[5117] + MEM[9825];
assign MEM[24041] = MEM[5122] + MEM[11702];
assign MEM[24042] = MEM[5125] + MEM[14141];
assign MEM[24043] = MEM[5140] + MEM[12367];
assign MEM[24044] = MEM[5142] + MEM[12368];
assign MEM[24045] = MEM[5151] + MEM[12580];
assign MEM[24046] = MEM[5167] + MEM[9755];
assign MEM[24047] = MEM[5173] + MEM[10057];
assign MEM[24048] = MEM[5178] + MEM[13866];
assign MEM[24049] = MEM[5191] + MEM[8647];
assign MEM[24050] = MEM[5197] + MEM[11773];
assign MEM[24051] = MEM[5198] + MEM[5914];
assign MEM[24052] = MEM[5202] + MEM[9092];
assign MEM[24053] = MEM[5207] + MEM[12126];
assign MEM[24054] = MEM[5212] + MEM[5736];
assign MEM[24055] = MEM[5219] + MEM[10456];
assign MEM[24056] = MEM[5228] + MEM[7656];
assign MEM[24057] = MEM[5245] + MEM[10659];
assign MEM[24058] = MEM[5259] + MEM[12715];
assign MEM[24059] = MEM[5269] + MEM[7107];
assign MEM[24060] = MEM[5284] + MEM[13770];
assign MEM[24061] = MEM[5293] + MEM[9714];
assign MEM[24062] = MEM[5298] + MEM[9207];
assign MEM[24063] = MEM[5299] + MEM[10410];
assign MEM[24064] = MEM[5301] + MEM[6189];
assign MEM[24065] = MEM[5302] + MEM[9817];
assign MEM[24066] = MEM[5304] + MEM[5470];
assign MEM[24067] = MEM[5311] + MEM[9537];
assign MEM[24068] = MEM[5312] + MEM[10510];
assign MEM[24069] = MEM[5315] + MEM[11778];
assign MEM[24070] = MEM[5326] + MEM[12389];
assign MEM[24071] = MEM[5330] + MEM[9206];
assign MEM[24072] = MEM[5339] + MEM[11634];
assign MEM[24073] = MEM[5347] + MEM[12331];
assign MEM[24074] = MEM[5354] + MEM[6419];
assign MEM[24075] = MEM[5381] + MEM[11109];
assign MEM[24076] = MEM[5390] + MEM[6094];
assign MEM[24077] = MEM[5399] + MEM[12319];
assign MEM[24078] = MEM[5404] + MEM[5516];
assign MEM[24079] = MEM[5405] + MEM[7443];
assign MEM[24080] = MEM[5426] + MEM[6078];
assign MEM[24081] = MEM[5439] + MEM[11847];
assign MEM[24082] = MEM[5443] + MEM[10853];
assign MEM[24083] = MEM[5446] + MEM[10643];
assign MEM[24084] = MEM[5451] + MEM[9798];
assign MEM[24085] = MEM[5452] + MEM[13074];
assign MEM[24086] = MEM[5461] + MEM[9331];
assign MEM[24087] = MEM[5469] + MEM[7167];
assign MEM[24088] = MEM[5474] + MEM[11851];
assign MEM[24089] = MEM[5479] + MEM[8766];
assign MEM[24090] = MEM[5483] + MEM[12485];
assign MEM[24091] = MEM[5499] + MEM[14898];
assign MEM[24092] = MEM[5500] + MEM[10370];
assign MEM[24093] = MEM[5511] + MEM[6858];
assign MEM[24094] = MEM[5523] + MEM[13058];
assign MEM[24095] = MEM[5524] + MEM[11239];
assign MEM[24096] = MEM[5526] + MEM[10839];
assign MEM[24097] = MEM[5530] + MEM[7085];
assign MEM[24098] = MEM[5540] + MEM[6111];
assign MEM[24099] = MEM[5549] + MEM[8873];
assign MEM[24100] = MEM[5555] + MEM[10537];
assign MEM[24101] = MEM[5571] + MEM[8318];
assign MEM[24102] = MEM[5580] + MEM[13277];
assign MEM[24103] = MEM[5606] + MEM[11588];
assign MEM[24104] = MEM[5614] + MEM[6753];
assign MEM[24105] = MEM[5615] + MEM[5990];
assign MEM[24106] = MEM[5621] + MEM[8273];
assign MEM[24107] = MEM[5623] + MEM[9855];
assign MEM[24108] = MEM[5634] + MEM[10071];
assign MEM[24109] = MEM[5635] + MEM[8497];
assign MEM[24110] = MEM[5641] + MEM[10055];
assign MEM[24111] = MEM[5642] + MEM[7849];
assign MEM[24112] = MEM[5650] + MEM[10470];
assign MEM[24113] = MEM[5652] + MEM[12322];
assign MEM[24114] = MEM[5658] + MEM[6904];
assign MEM[24115] = MEM[5659] + MEM[6343];
assign MEM[24116] = MEM[5666] + MEM[7871];
assign MEM[24117] = MEM[5669] + MEM[8723];
assign MEM[24118] = MEM[5674] + MEM[5782];
assign MEM[24119] = MEM[5684] + MEM[7529];
assign MEM[24120] = MEM[5692] + MEM[11687];
assign MEM[24121] = MEM[5694] + MEM[12259];
assign MEM[24122] = MEM[5698] + MEM[6307];
assign MEM[24123] = MEM[5702] + MEM[8977];
assign MEM[24124] = MEM[5703] + MEM[8533];
assign MEM[24125] = MEM[5711] + MEM[6031];
assign MEM[24126] = MEM[5747] + MEM[10861];
assign MEM[24127] = MEM[5754] + MEM[11173];
assign MEM[24128] = MEM[5756] + MEM[12244];
assign MEM[24129] = MEM[5763] + MEM[11558];
assign MEM[24130] = MEM[5766] + MEM[8389];
assign MEM[24131] = MEM[5774] + MEM[13390];
assign MEM[24132] = MEM[5780] + MEM[12239];
assign MEM[24133] = MEM[5786] + MEM[10207];
assign MEM[24134] = MEM[5794] + MEM[6723];
assign MEM[24135] = MEM[5807] + MEM[8513];
assign MEM[24136] = MEM[5845] + MEM[8913];
assign MEM[24137] = MEM[5846] + MEM[6279];
assign MEM[24138] = MEM[5847] + MEM[7043];
assign MEM[24139] = MEM[5861] + MEM[9911];
assign MEM[24140] = MEM[5862] + MEM[6784];
assign MEM[24141] = MEM[5875] + MEM[13679];
assign MEM[24142] = MEM[5899] + MEM[7707];
assign MEM[24143] = MEM[5901] + MEM[11939];
assign MEM[24144] = MEM[5904] + MEM[6703];
assign MEM[24145] = MEM[5911] + MEM[7050];
assign MEM[24146] = MEM[5923] + MEM[16156];
assign MEM[24147] = MEM[5934] + MEM[13225];
assign MEM[24148] = MEM[5936] + MEM[7448];
assign MEM[24149] = MEM[5937] + MEM[10006];
assign MEM[24150] = MEM[5938] + MEM[6336];
assign MEM[24151] = MEM[5943] + MEM[6298];
assign MEM[24152] = MEM[5946] + MEM[6425];
assign MEM[24153] = MEM[5949] + MEM[13160];
assign MEM[24154] = MEM[5952] + MEM[6556];
assign MEM[24155] = MEM[5956] + MEM[13405];
assign MEM[24156] = MEM[5962] + MEM[6888];
assign MEM[24157] = MEM[5963] + MEM[12318];
assign MEM[24158] = MEM[5970] + MEM[13844];
assign MEM[24159] = MEM[5973] + MEM[11007];
assign MEM[24160] = MEM[5981] + MEM[10414];
assign MEM[24161] = MEM[5986] + MEM[13125];
assign MEM[24162] = MEM[5989] + MEM[12932];
assign MEM[24163] = MEM[6005] + MEM[12250];
assign MEM[24164] = MEM[6011] + MEM[9321];
assign MEM[24165] = MEM[6014] + MEM[9934];
assign MEM[24166] = MEM[6045] + MEM[6487];
assign MEM[24167] = MEM[6046] + MEM[11053];
assign MEM[24168] = MEM[6047] + MEM[6598];
assign MEM[24169] = MEM[6077] + MEM[10560];
assign MEM[24170] = MEM[6087] + MEM[6473];
assign MEM[24171] = MEM[6102] + MEM[7343];
assign MEM[24172] = MEM[6115] + MEM[10670];
assign MEM[24173] = MEM[6119] + MEM[10473];
assign MEM[24174] = MEM[6123] + MEM[6272];
assign MEM[24175] = MEM[6125] + MEM[14336];
assign MEM[24176] = MEM[6127] + MEM[11541];
assign MEM[24177] = MEM[6130] + MEM[14082];
assign MEM[24178] = MEM[6135] + MEM[9125];
assign MEM[24179] = MEM[6141] + MEM[10467];
assign MEM[24180] = MEM[6147] + MEM[7663];
assign MEM[24181] = MEM[6149] + MEM[11655];
assign MEM[24182] = MEM[6157] + MEM[11187];
assign MEM[24183] = MEM[6163] + MEM[11991];
assign MEM[24184] = MEM[6165] + MEM[9756];
assign MEM[24185] = MEM[6166] + MEM[13489];
assign MEM[24186] = MEM[6167] + MEM[8641];
assign MEM[24187] = MEM[6170] + MEM[6964];
assign MEM[24188] = MEM[6171] + MEM[14493];
assign MEM[24189] = MEM[6174] + MEM[9878];
assign MEM[24190] = MEM[6175] + MEM[11797];
assign MEM[24191] = MEM[6181] + MEM[7797];
assign MEM[24192] = MEM[6182] + MEM[6877];
assign MEM[24193] = MEM[6188] + MEM[13352];
assign MEM[24194] = MEM[6191] + MEM[7057];
assign MEM[24195] = MEM[6195] + MEM[10619];
assign MEM[24196] = MEM[6198] + MEM[6415];
assign MEM[24197] = MEM[6203] + MEM[10557];
assign MEM[24198] = MEM[6214] + MEM[9194];
assign MEM[24199] = MEM[6215] + MEM[10776];
assign MEM[24200] = MEM[6219] + MEM[6582];
assign MEM[24201] = MEM[6220] + MEM[7316];
assign MEM[24202] = MEM[6228] + MEM[9294];
assign MEM[24203] = MEM[6237] + MEM[10608];
assign MEM[24204] = MEM[6238] + MEM[8229];
assign MEM[24205] = MEM[6239] + MEM[11994];
assign MEM[24206] = MEM[6253] + MEM[7562];
assign MEM[24207] = MEM[6261] + MEM[12359];
assign MEM[24208] = MEM[6262] + MEM[10589];
assign MEM[24209] = MEM[6274] + MEM[9081];
assign MEM[24210] = MEM[6291] + MEM[7841];
assign MEM[24211] = MEM[6305] + MEM[7559];
assign MEM[24212] = MEM[6308] + MEM[9806];
assign MEM[24213] = MEM[6317] + MEM[6462];
assign MEM[24214] = MEM[6324] + MEM[13498];
assign MEM[24215] = MEM[6329] + MEM[10750];
assign MEM[24216] = MEM[6330] + MEM[8365];
assign MEM[24217] = MEM[6371] + MEM[8930];
assign MEM[24218] = MEM[6372] + MEM[10099];
assign MEM[24219] = MEM[6381] + MEM[13755];
assign MEM[24220] = MEM[6391] + MEM[11673];
assign MEM[24221] = MEM[6416] + MEM[12222];
assign MEM[24222] = MEM[6421] + MEM[11706];
assign MEM[24223] = MEM[6429] + MEM[7279];
assign MEM[24224] = MEM[6431] + MEM[12269];
assign MEM[24225] = MEM[6434] + MEM[11015];
assign MEM[24226] = MEM[6438] + MEM[10246];
assign MEM[24227] = MEM[6439] + MEM[11979];
assign MEM[24228] = MEM[6442] + MEM[13466];
assign MEM[24229] = MEM[6443] + MEM[9195];
assign MEM[24230] = MEM[6453] + MEM[12758];
assign MEM[24231] = MEM[6466] + MEM[11643];
assign MEM[24232] = MEM[6485] + MEM[10620];
assign MEM[24233] = MEM[6513] + MEM[10430];
assign MEM[24234] = MEM[6518] + MEM[12138];
assign MEM[24235] = MEM[6532] + MEM[6843];
assign MEM[24236] = MEM[6555] + MEM[11192];
assign MEM[24237] = MEM[6560] + MEM[10983];
assign MEM[24238] = MEM[6562] + MEM[10876];
assign MEM[24239] = MEM[6566] + MEM[13159];
assign MEM[24240] = MEM[6580] + MEM[7090];
assign MEM[24241] = MEM[6586] + MEM[12394];
assign MEM[24242] = MEM[6587] + MEM[7319];
assign MEM[24243] = MEM[6593] + MEM[6902];
assign MEM[24244] = MEM[6597] + MEM[10300];
assign MEM[24245] = MEM[6610] + MEM[10069];
assign MEM[24246] = MEM[6611] + MEM[10667];
assign MEM[24247] = MEM[6618] + MEM[7012];
assign MEM[24248] = MEM[6634] + MEM[10381];
assign MEM[24249] = MEM[6648] + MEM[10519];
assign MEM[24250] = MEM[6650] + MEM[10366];
assign MEM[24251] = MEM[6652] + MEM[15107];
assign MEM[24252] = MEM[6656] + MEM[11697];
assign MEM[24253] = MEM[6667] + MEM[10844];
assign MEM[24254] = MEM[6670] + MEM[6846];
assign MEM[24255] = MEM[6671] + MEM[8523];
assign MEM[24256] = MEM[6674] + MEM[12850];
assign MEM[24257] = MEM[6676] + MEM[8325];
assign MEM[24258] = MEM[6683] + MEM[10716];
assign MEM[24259] = MEM[6684] + MEM[8274];
assign MEM[24260] = MEM[6691] + MEM[10636];
assign MEM[24261] = MEM[6698] + MEM[8615];
assign MEM[24262] = MEM[6699] + MEM[7395];
assign MEM[24263] = MEM[6700] + MEM[11383];
assign MEM[24264] = MEM[6710] + MEM[10336];
assign MEM[24265] = MEM[6715] + MEM[10367];
assign MEM[24266] = MEM[6717] + MEM[7384];
assign MEM[24267] = MEM[6722] + MEM[7517];
assign MEM[24268] = MEM[6736] + MEM[10490];
assign MEM[24269] = MEM[6744] + MEM[9576];
assign MEM[24270] = MEM[6745] + MEM[12397];
assign MEM[24271] = MEM[6751] + MEM[6956];
assign MEM[24272] = MEM[6754] + MEM[13032];
assign MEM[24273] = MEM[6755] + MEM[10453];
assign MEM[24274] = MEM[6776] + MEM[15899];
assign MEM[24275] = MEM[6778] + MEM[8431];
assign MEM[24276] = MEM[6785] + MEM[8652];
assign MEM[24277] = MEM[6801] + MEM[8604];
assign MEM[24278] = MEM[6805] + MEM[11483];
assign MEM[24279] = MEM[6810] + MEM[10409];
assign MEM[24280] = MEM[6818] + MEM[17198];
assign MEM[24281] = MEM[6823] + MEM[8183];
assign MEM[24282] = MEM[6829] + MEM[7728];
assign MEM[24283] = MEM[6837] + MEM[15761];
assign MEM[24284] = MEM[6841] + MEM[8079];
assign MEM[24285] = MEM[6842] + MEM[7645];
assign MEM[24286] = MEM[6847] + MEM[7086];
assign MEM[24287] = MEM[6848] + MEM[6982];
assign MEM[24288] = MEM[6853] + MEM[13760];
assign MEM[24289] = MEM[6855] + MEM[10584];
assign MEM[24290] = MEM[6858] + MEM[16240];
assign MEM[24291] = MEM[6864] + MEM[7236];
assign MEM[24292] = MEM[6875] + MEM[8440];
assign MEM[24293] = MEM[6878] + MEM[9000];
assign MEM[24294] = MEM[6881] + MEM[10032];
assign MEM[24295] = MEM[6893] + MEM[9869];
assign MEM[24296] = MEM[6907] + MEM[8267];
assign MEM[24297] = MEM[6910] + MEM[10536];
assign MEM[24298] = MEM[6923] + MEM[10058];
assign MEM[24299] = MEM[6929] + MEM[8598];
assign MEM[24300] = MEM[6938] + MEM[7092];
assign MEM[24301] = MEM[6941] + MEM[10913];
assign MEM[24302] = MEM[6945] + MEM[10347];
assign MEM[24303] = MEM[6953] + MEM[9827];
assign MEM[24304] = MEM[6962] + MEM[14928];
assign MEM[24305] = MEM[6963] + MEM[7859];
assign MEM[24306] = MEM[6967] + MEM[7440];
assign MEM[24307] = MEM[6968] + MEM[14100];
assign MEM[24308] = MEM[6969] + MEM[9453];
assign MEM[24309] = MEM[6974] + MEM[12509];
assign MEM[24310] = MEM[6981] + MEM[7890];
assign MEM[24311] = MEM[6993] + MEM[7060];
assign MEM[24312] = MEM[6999] + MEM[12349];
assign MEM[24313] = MEM[7000] + MEM[12084];
assign MEM[24314] = MEM[7003] + MEM[13279];
assign MEM[24315] = MEM[7011] + MEM[11791];
assign MEM[24316] = MEM[7017] + MEM[11157];
assign MEM[24317] = MEM[7029] + MEM[7945];
assign MEM[24318] = MEM[7031] + MEM[9723];
assign MEM[24319] = MEM[7032] + MEM[9955];
assign MEM[24320] = MEM[7044] + MEM[12482];
assign MEM[24321] = MEM[7047] + MEM[11124];
assign MEM[24322] = MEM[7061] + MEM[7456];
assign MEM[24323] = MEM[7063] + MEM[9287];
assign MEM[24324] = MEM[7070] + MEM[11551];
assign MEM[24325] = MEM[7071] + MEM[12446];
assign MEM[24326] = MEM[7088] + MEM[8754];
assign MEM[24327] = MEM[7095] + MEM[11125];
assign MEM[24328] = MEM[7096] + MEM[9829];
assign MEM[24329] = MEM[7103] + MEM[17702];
assign MEM[24330] = MEM[7119] + MEM[7248];
assign MEM[24331] = MEM[7121] + MEM[7595];
assign MEM[24332] = MEM[7124] + MEM[11354];
assign MEM[24333] = MEM[7125] + MEM[16741];
assign MEM[24334] = MEM[7143] + MEM[7978];
assign MEM[24335] = MEM[7145] + MEM[8294];
assign MEM[24336] = MEM[7146] + MEM[13447];
assign MEM[24337] = MEM[7148] + MEM[7743];
assign MEM[24338] = MEM[7150] + MEM[9062];
assign MEM[24339] = MEM[7152] + MEM[8535];
assign MEM[24340] = MEM[7154] + MEM[8090];
assign MEM[24341] = MEM[7166] + MEM[8650];
assign MEM[24342] = MEM[7173] + MEM[9053];
assign MEM[24343] = MEM[7197] + MEM[15715];
assign MEM[24344] = MEM[7198] + MEM[7233];
assign MEM[24345] = MEM[7203] + MEM[10932];
assign MEM[24346] = MEM[7204] + MEM[10045];
assign MEM[24347] = MEM[7205] + MEM[8324];
assign MEM[24348] = MEM[7207] + MEM[14216];
assign MEM[24349] = MEM[7210] + MEM[15886];
assign MEM[24350] = MEM[7214] + MEM[13134];
assign MEM[24351] = MEM[7215] + MEM[13385];
assign MEM[24352] = MEM[7238] + MEM[12062];
assign MEM[24353] = MEM[7240] + MEM[12518];
assign MEM[24354] = MEM[7245] + MEM[10884];
assign MEM[24355] = MEM[7250] + MEM[13221];
assign MEM[24356] = MEM[7255] + MEM[10588];
assign MEM[24357] = MEM[7256] + MEM[9327];
assign MEM[24358] = MEM[7273] + MEM[11668];
assign MEM[24359] = MEM[7283] + MEM[12408];
assign MEM[24360] = MEM[7294] + MEM[11219];
assign MEM[24361] = MEM[7295] + MEM[12298];
assign MEM[24362] = MEM[7298] + MEM[8248];
assign MEM[24363] = MEM[7303] + MEM[11375];
assign MEM[24364] = MEM[7315] + MEM[8992];
assign MEM[24365] = MEM[7320] + MEM[10005];
assign MEM[24366] = MEM[7326] + MEM[9499];
assign MEM[24367] = MEM[7327] + MEM[9463];
assign MEM[24368] = MEM[7330] + MEM[12528];
assign MEM[24369] = MEM[7334] + MEM[10021];
assign MEM[24370] = MEM[7350] + MEM[12060];
assign MEM[24371] = MEM[7353] + MEM[11070];
assign MEM[24372] = MEM[7355] + MEM[9761];
assign MEM[24373] = MEM[7359] + MEM[8006];
assign MEM[24374] = MEM[7364] + MEM[15735];
assign MEM[24375] = MEM[7365] + MEM[8949];
assign MEM[24376] = MEM[7367] + MEM[11408];
assign MEM[24377] = MEM[7376] + MEM[11982];
assign MEM[24378] = MEM[7377] + MEM[11009];
assign MEM[24379] = MEM[7378] + MEM[10403];
assign MEM[24380] = MEM[7379] + MEM[13394];
assign MEM[24381] = MEM[7387] + MEM[13520];
assign MEM[24382] = MEM[7389] + MEM[13112];
assign MEM[24383] = MEM[7394] + MEM[9104];
assign MEM[24384] = MEM[7407] + MEM[12500];
assign MEM[24385] = MEM[7418] + MEM[12007];
assign MEM[24386] = MEM[7419] + MEM[9376];
assign MEM[24387] = MEM[7421] + MEM[17699];
assign MEM[24388] = MEM[7424] + MEM[13476];
assign MEM[24389] = MEM[7431] + MEM[12708];
assign MEM[24390] = MEM[7434] + MEM[8101];
assign MEM[24391] = MEM[7436] + MEM[9736];
assign MEM[24392] = MEM[7446] + MEM[8226];
assign MEM[24393] = MEM[7449] + MEM[11145];
assign MEM[24394] = MEM[7453] + MEM[10152];
assign MEM[24395] = MEM[7458] + MEM[9372];
assign MEM[24396] = MEM[7465] + MEM[12400];
assign MEM[24397] = MEM[7467] + MEM[14245];
assign MEM[24398] = MEM[7468] + MEM[9311];
assign MEM[24399] = MEM[7484] + MEM[8529];
assign MEM[24400] = MEM[7485] + MEM[8960];
assign MEM[24401] = MEM[7504] + MEM[9612];
assign MEM[24402] = MEM[7505] + MEM[7994];
assign MEM[24403] = MEM[7519] + MEM[9938];
assign MEM[24404] = MEM[7524] + MEM[12619];
assign MEM[24405] = MEM[7535] + MEM[11142];
assign MEM[24406] = MEM[7551] + MEM[12748];
assign MEM[24407] = MEM[7560] + MEM[9201];
assign MEM[24408] = MEM[7568] + MEM[12693];
assign MEM[24409] = MEM[7569] + MEM[9817];
assign MEM[24410] = MEM[7572] + MEM[10131];
assign MEM[24411] = MEM[7578] + MEM[11973];
assign MEM[24412] = MEM[7579] + MEM[14286];
assign MEM[24413] = MEM[7600] + MEM[12247];
assign MEM[24414] = MEM[7601] + MEM[9472];
assign MEM[24415] = MEM[7603] + MEM[8520];
assign MEM[24416] = MEM[7608] + MEM[8118];
assign MEM[24417] = MEM[7609] + MEM[10770];
assign MEM[24418] = MEM[7616] + MEM[10664];
assign MEM[24419] = MEM[7618] + MEM[15394];
assign MEM[24420] = MEM[7628] + MEM[11151];
assign MEM[24421] = MEM[7629] + MEM[11961];
assign MEM[24422] = MEM[7633] + MEM[12080];
assign MEM[24423] = MEM[7655] + MEM[11516];
assign MEM[24424] = MEM[7662] + MEM[8170];
assign MEM[24425] = MEM[7663] + MEM[10909];
assign MEM[24426] = MEM[7675] + MEM[12927];
assign MEM[24427] = MEM[7678] + MEM[9206];
assign MEM[24428] = MEM[7679] + MEM[10376];
assign MEM[24429] = MEM[7680] + MEM[12292];
assign MEM[24430] = MEM[7687] + MEM[13272];
assign MEM[24431] = MEM[7694] + MEM[9400];
assign MEM[24432] = MEM[7697] + MEM[9585];
assign MEM[24433] = MEM[7699] + MEM[10723];
assign MEM[24434] = MEM[7705] + MEM[10936];
assign MEM[24435] = MEM[7712] + MEM[13301];
assign MEM[24436] = MEM[7714] + MEM[12853];
assign MEM[24437] = MEM[7715] + MEM[10464];
assign MEM[24438] = MEM[7716] + MEM[12838];
assign MEM[24439] = MEM[7723] + MEM[9055];
assign MEM[24440] = MEM[7725] + MEM[13176];
assign MEM[24441] = MEM[7726] + MEM[13954];
assign MEM[24442] = MEM[7732] + MEM[11047];
assign MEM[24443] = MEM[7734] + MEM[8178];
assign MEM[24444] = MEM[7737] + MEM[7933];
assign MEM[24445] = MEM[7747] + MEM[11431];
assign MEM[24446] = MEM[7748] + MEM[13164];
assign MEM[24447] = MEM[7750] + MEM[8132];
assign MEM[24448] = MEM[7754] + MEM[9439];
assign MEM[24449] = MEM[7755] + MEM[15931];
assign MEM[24450] = MEM[7761] + MEM[9910];
assign MEM[24451] = MEM[7766] + MEM[11049];
assign MEM[24452] = MEM[7769] + MEM[13572];
assign MEM[24453] = MEM[7770] + MEM[11929];
assign MEM[24454] = MEM[7779] + MEM[12652];
assign MEM[24455] = MEM[7793] + MEM[8811];
assign MEM[24456] = MEM[7801] + MEM[11076];
assign MEM[24457] = MEM[7837] + MEM[16286];
assign MEM[24458] = MEM[7840] + MEM[13154];
assign MEM[24459] = MEM[7845] + MEM[10404];
assign MEM[24460] = MEM[7847] + MEM[7956];
assign MEM[24461] = MEM[7848] + MEM[12689];
assign MEM[24462] = MEM[7856] + MEM[11943];
assign MEM[24463] = MEM[7863] + MEM[16087];
assign MEM[24464] = MEM[7865] + MEM[8691];
assign MEM[24465] = MEM[7867] + MEM[10358];
assign MEM[24466] = MEM[7880] + MEM[9038];
assign MEM[24467] = MEM[7888] + MEM[13706];
assign MEM[24468] = MEM[7908] + MEM[10902];
assign MEM[24469] = MEM[7909] + MEM[8311];
assign MEM[24470] = MEM[7910] + MEM[8889];
assign MEM[24471] = MEM[7927] + MEM[9995];
assign MEM[24472] = MEM[7937] + MEM[9796];
assign MEM[24473] = MEM[7949] + MEM[12718];
assign MEM[24474] = MEM[7965] + MEM[8285];
assign MEM[24475] = MEM[7972] + MEM[13756];
assign MEM[24476] = MEM[7973] + MEM[12337];
assign MEM[24477] = MEM[7985] + MEM[8750];
assign MEM[24478] = MEM[7987] + MEM[12701];
assign MEM[24479] = MEM[7988] + MEM[11310];
assign MEM[24480] = MEM[7993] + MEM[11981];
assign MEM[24481] = MEM[7998] + MEM[10823];
assign MEM[24482] = MEM[8001] + MEM[10399];
assign MEM[24483] = MEM[8002] + MEM[10998];
assign MEM[24484] = MEM[8007] + MEM[8280];
assign MEM[24485] = MEM[8009] + MEM[10757];
assign MEM[24486] = MEM[8013] + MEM[9399];
assign MEM[24487] = MEM[8014] + MEM[8023];
assign MEM[24488] = MEM[8016] + MEM[8425];
assign MEM[24489] = MEM[8018] + MEM[9326];
assign MEM[24490] = MEM[8022] + MEM[10556];
assign MEM[24491] = MEM[8028] + MEM[11754];
assign MEM[24492] = MEM[8029] + MEM[10223];
assign MEM[24493] = MEM[8036] + MEM[13456];
assign MEM[24494] = MEM[8040] + MEM[10369];
assign MEM[24495] = MEM[8041] + MEM[15036];
assign MEM[24496] = MEM[8046] + MEM[12401];
assign MEM[24497] = MEM[8048] + MEM[11137];
assign MEM[24498] = MEM[8051] + MEM[12370];
assign MEM[24499] = MEM[8059] + MEM[11328];
assign MEM[24500] = MEM[8063] + MEM[11001];
assign MEM[24501] = MEM[8071] + MEM[9811];
assign MEM[24502] = MEM[8072] + MEM[10468];
assign MEM[24503] = MEM[8073] + MEM[13686];
assign MEM[24504] = MEM[8075] + MEM[11955];
assign MEM[24505] = MEM[8080] + MEM[12113];
assign MEM[24506] = MEM[8084] + MEM[10692];
assign MEM[24507] = MEM[8095] + MEM[11302];
assign MEM[24508] = MEM[8103] + MEM[12046];
assign MEM[24509] = MEM[8110] + MEM[10406];
assign MEM[24510] = MEM[8122] + MEM[8147];
assign MEM[24511] = MEM[8125] + MEM[15174];
assign MEM[24512] = MEM[8130] + MEM[9049];
assign MEM[24513] = MEM[8134] + MEM[10896];
assign MEM[24514] = MEM[8136] + MEM[9767];
assign MEM[24515] = MEM[8142] + MEM[10579];
assign MEM[24516] = MEM[8143] + MEM[12550];
assign MEM[24517] = MEM[8145] + MEM[10959];
assign MEM[24518] = MEM[8155] + MEM[11465];
assign MEM[24519] = MEM[8164] + MEM[12945];
assign MEM[24520] = MEM[8169] + MEM[11874];
assign MEM[24521] = MEM[8177] + MEM[11422];
assign MEM[24522] = MEM[8181] + MEM[10278];
assign MEM[24523] = MEM[8184] + MEM[8620];
assign MEM[24524] = MEM[8186] + MEM[8743];
assign MEM[24525] = MEM[8187] + MEM[14019];
assign MEM[24526] = MEM[8193] + MEM[8348];
assign MEM[24527] = MEM[8194] + MEM[10618];
assign MEM[24528] = MEM[8200] + MEM[9054];
assign MEM[24529] = MEM[8201] + MEM[8643];
assign MEM[24530] = MEM[8202] + MEM[10465];
assign MEM[24531] = MEM[8204] + MEM[13748];
assign MEM[24532] = MEM[8207] + MEM[10869];
assign MEM[24533] = MEM[8210] + MEM[10102];
assign MEM[24534] = MEM[8211] + MEM[12794];
assign MEM[24535] = MEM[8213] + MEM[13587];
assign MEM[24536] = MEM[8215] + MEM[11601];
assign MEM[24537] = MEM[8216] + MEM[12732];
assign MEM[24538] = MEM[8233] + MEM[8581];
assign MEM[24539] = MEM[8233] + MEM[10754];
assign MEM[24540] = MEM[8238] + MEM[10386];
assign MEM[24541] = MEM[8240] + MEM[13189];
assign MEM[24542] = MEM[8252] + MEM[10782];
assign MEM[24543] = MEM[8255] + MEM[10801];
assign MEM[24544] = MEM[8257] + MEM[10433];
assign MEM[24545] = MEM[8261] + MEM[11724];
assign MEM[24546] = MEM[8271] + MEM[10482];
assign MEM[24547] = MEM[8272] + MEM[11618];
assign MEM[24548] = MEM[8278] + MEM[13015];
assign MEM[24549] = MEM[8279] + MEM[11887];
assign MEM[24550] = MEM[8292] + MEM[8499];
assign MEM[24551] = MEM[8298] + MEM[10177];
assign MEM[24552] = MEM[8302] + MEM[11631];
assign MEM[24553] = MEM[8322] + MEM[10097];
assign MEM[24554] = MEM[8334] + MEM[10805];
assign MEM[24555] = MEM[8356] + MEM[12578];
assign MEM[24556] = MEM[8359] + MEM[11671];
assign MEM[24557] = MEM[8360] + MEM[10276];
assign MEM[24558] = MEM[8376] + MEM[11548];
assign MEM[24559] = MEM[8377] + MEM[10440];
assign MEM[24560] = MEM[8396] + MEM[10915];
assign MEM[24561] = MEM[8411] + MEM[9147];
assign MEM[24562] = MEM[8414] + MEM[16046];
assign MEM[24563] = MEM[8416] + MEM[15521];
assign MEM[24564] = MEM[8418] + MEM[11808];
assign MEM[24565] = MEM[8428] + MEM[13064];
assign MEM[24566] = MEM[8439] + MEM[13004];
assign MEM[24567] = MEM[8442] + MEM[10944];
assign MEM[24568] = MEM[8457] + MEM[16339];
assign MEM[24569] = MEM[8465] + MEM[8820];
assign MEM[24570] = MEM[8466] + MEM[11966];
assign MEM[24571] = MEM[8467] + MEM[11868];
assign MEM[24572] = MEM[8469] + MEM[11800];
assign MEM[24573] = MEM[8473] + MEM[8498];
assign MEM[24574] = MEM[8474] + MEM[9732];
assign MEM[24575] = MEM[8476] + MEM[14298];
assign MEM[24576] = MEM[8490] + MEM[15756];
assign MEM[24577] = MEM[8492] + MEM[10327];
assign MEM[24578] = MEM[8493] + MEM[12879];
assign MEM[24579] = MEM[8499] + MEM[13404];
assign MEM[24580] = MEM[8503] + MEM[11309];
assign MEM[24581] = MEM[8510] + MEM[9130];
assign MEM[24582] = MEM[8510] + MEM[12999];
assign MEM[24583] = MEM[8514] + MEM[16104];
assign MEM[24584] = MEM[8516] + MEM[14503];
assign MEM[24585] = MEM[8517] + MEM[12069];
assign MEM[24586] = MEM[8545] + MEM[8860];
assign MEM[24587] = MEM[8551] + MEM[9595];
assign MEM[24588] = MEM[8552] + MEM[13135];
assign MEM[24589] = MEM[8557] + MEM[12364];
assign MEM[24590] = MEM[8558] + MEM[12634];
assign MEM[24591] = MEM[8560] + MEM[12163];
assign MEM[24592] = MEM[8565] + MEM[10758];
assign MEM[24593] = MEM[8571] + MEM[8886];
assign MEM[24594] = MEM[8572] + MEM[10705];
assign MEM[24595] = MEM[8574] + MEM[10892];
assign MEM[24596] = MEM[8576] + MEM[10481];
assign MEM[24597] = MEM[8586] + MEM[10273];
assign MEM[24598] = MEM[8587] + MEM[12152];
assign MEM[24599] = MEM[8600] + MEM[10634];
assign MEM[24600] = MEM[8602] + MEM[15203];
assign MEM[24601] = MEM[8608] + MEM[8632];
assign MEM[24602] = MEM[8612] + MEM[9417];
assign MEM[24603] = MEM[8613] + MEM[13446];
assign MEM[24604] = MEM[8614] + MEM[10077];
assign MEM[24605] = MEM[8618] + MEM[14315];
assign MEM[24606] = MEM[8621] + MEM[11822];
assign MEM[24607] = MEM[8626] + MEM[9722];
assign MEM[24608] = MEM[8631] + MEM[10663];
assign MEM[24609] = MEM[8636] + MEM[11080];
assign MEM[24610] = MEM[8637] + MEM[10136];
assign MEM[24611] = MEM[8648] + MEM[12682];
assign MEM[24612] = MEM[8649] + MEM[12878];
assign MEM[24613] = MEM[8654] + MEM[12199];
assign MEM[24614] = MEM[8671] + MEM[9173];
assign MEM[24615] = MEM[8673] + MEM[10321];
assign MEM[24616] = MEM[8675] + MEM[8835];
assign MEM[24617] = MEM[8692] + MEM[10674];
assign MEM[24618] = MEM[8693] + MEM[12752];
assign MEM[24619] = MEM[8709] + MEM[11882];
assign MEM[24620] = MEM[8712] + MEM[9754];
assign MEM[24621] = MEM[8734] + MEM[13753];
assign MEM[24622] = MEM[8735] + MEM[9966];
assign MEM[24623] = MEM[8737] + MEM[15067];
assign MEM[24624] = MEM[8739] + MEM[8890];
assign MEM[24625] = MEM[8739] + MEM[17370];
assign MEM[24626] = MEM[8746] + MEM[8950];
assign MEM[24627] = MEM[8759] + MEM[11263];
assign MEM[24628] = MEM[8762] + MEM[12937];
assign MEM[24629] = MEM[8763] + MEM[12148];
assign MEM[24630] = MEM[8767] + MEM[12079];
assign MEM[24631] = MEM[8770] + MEM[14622];
assign MEM[24632] = MEM[8772] + MEM[8861];
assign MEM[24633] = MEM[8774] + MEM[12450];
assign MEM[24634] = MEM[8778] + MEM[9912];
assign MEM[24635] = MEM[8795] + MEM[10845];
assign MEM[24636] = MEM[8801] + MEM[9784];
assign MEM[24637] = MEM[8802] + MEM[14738];
assign MEM[24638] = MEM[8818] + MEM[10581];
assign MEM[24639] = MEM[8827] + MEM[10673];
assign MEM[24640] = MEM[8830] + MEM[10353];
assign MEM[24641] = MEM[8833] + MEM[12288];
assign MEM[24642] = MEM[8841] + MEM[13823];
assign MEM[24643] = MEM[8842] + MEM[16911];
assign MEM[24644] = MEM[8844] + MEM[12184];
assign MEM[24645] = MEM[8848] + MEM[11638];
assign MEM[24646] = MEM[8853] + MEM[11853];
assign MEM[24647] = MEM[8854] + MEM[10295];
assign MEM[24648] = MEM[8858] + MEM[12714];
assign MEM[24649] = MEM[8864] + MEM[10222];
assign MEM[24650] = MEM[8874] + MEM[10485];
assign MEM[24651] = MEM[8882] + MEM[11067];
assign MEM[24652] = MEM[8887] + MEM[15363];
assign MEM[24653] = MEM[8888] + MEM[10229];
assign MEM[24654] = MEM[8891] + MEM[12022];
assign MEM[24655] = MEM[8892] + MEM[11129];
assign MEM[24656] = MEM[8901] + MEM[11856];
assign MEM[24657] = MEM[8904] + MEM[9874];
assign MEM[24658] = MEM[8906] + MEM[12495];
assign MEM[24659] = MEM[8915] + MEM[9149];
assign MEM[24660] = MEM[8925] + MEM[12562];
assign MEM[24661] = MEM[8928] + MEM[10443];
assign MEM[24662] = MEM[8928] + MEM[13899];
assign MEM[24663] = MEM[8929] + MEM[11713];
assign MEM[24664] = MEM[8934] + MEM[10022];
assign MEM[24665] = MEM[8940] + MEM[10524];
assign MEM[24666] = MEM[8955] + MEM[9654];
assign MEM[24667] = MEM[8960] + MEM[12033];
assign MEM[24668] = MEM[8961] + MEM[10339];
assign MEM[24669] = MEM[8973] + MEM[10322];
assign MEM[24670] = MEM[8986] + MEM[11220];
assign MEM[24671] = MEM[8994] + MEM[14538];
assign MEM[24672] = MEM[8995] + MEM[10860];
assign MEM[24673] = MEM[9006] + MEM[12162];
assign MEM[24674] = MEM[9008] + MEM[9320];
assign MEM[24675] = MEM[9015] + MEM[11176];
assign MEM[24676] = MEM[9022] + MEM[11013];
assign MEM[24677] = MEM[9023] + MEM[10918];
assign MEM[24678] = MEM[9037] + MEM[10281];
assign MEM[24679] = MEM[9041] + MEM[10952];
assign MEM[24680] = MEM[9045] + MEM[10749];
assign MEM[24681] = MEM[9058] + MEM[10831];
assign MEM[24682] = MEM[9068] + MEM[10038];
assign MEM[24683] = MEM[9069] + MEM[12309];
assign MEM[24684] = MEM[9080] + MEM[12216];
assign MEM[24685] = MEM[9087] + MEM[9964];
assign MEM[24686] = MEM[9088] + MEM[13699];
assign MEM[24687] = MEM[9103] + MEM[11880];
assign MEM[24688] = MEM[9110] + MEM[9843];
assign MEM[24689] = MEM[9120] + MEM[9166];
assign MEM[24690] = MEM[9139] + MEM[10743];
assign MEM[24691] = MEM[9142] + MEM[11663];
assign MEM[24692] = MEM[9145] + MEM[10418];
assign MEM[24693] = MEM[9157] + MEM[9483];
assign MEM[24694] = MEM[9165] + MEM[11204];
assign MEM[24695] = MEM[9169] + MEM[12506];
assign MEM[24696] = MEM[9175] + MEM[11917];
assign MEM[24697] = MEM[9183] + MEM[10836];
assign MEM[24698] = MEM[9184] + MEM[10759];
assign MEM[24699] = MEM[9185] + MEM[10239];
assign MEM[24700] = MEM[9187] + MEM[14042];
assign MEM[24701] = MEM[9204] + MEM[10677];
assign MEM[24702] = MEM[9208] + MEM[11225];
assign MEM[24703] = MEM[9210] + MEM[12303];
assign MEM[24704] = MEM[9212] + MEM[10865];
assign MEM[24705] = MEM[9231] + MEM[11024];
assign MEM[24706] = MEM[9243] + MEM[11133];
assign MEM[24707] = MEM[9248] + MEM[9257];
assign MEM[24708] = MEM[9258] + MEM[10644];
assign MEM[24709] = MEM[9277] + MEM[12235];
assign MEM[24710] = MEM[9278] + MEM[13897];
assign MEM[24711] = MEM[9299] + MEM[12414];
assign MEM[24712] = MEM[9310] + MEM[10695];
assign MEM[24713] = MEM[9317] + MEM[15141];
assign MEM[24714] = MEM[9330] + MEM[11253];
assign MEM[24715] = MEM[9331] + MEM[10833];
assign MEM[24716] = MEM[9344] + MEM[9908];
assign MEM[24717] = MEM[9346] + MEM[12694];
assign MEM[24718] = MEM[9350] + MEM[10031];
assign MEM[24719] = MEM[9354] + MEM[9632];
assign MEM[24720] = MEM[9370] + MEM[11050];
assign MEM[24721] = MEM[9373] + MEM[9518];
assign MEM[24722] = MEM[9384] + MEM[10478];
assign MEM[24723] = MEM[9388] + MEM[10953];
assign MEM[24724] = MEM[9406] + MEM[12228];
assign MEM[24725] = MEM[9407] + MEM[15207];
assign MEM[24726] = MEM[9416] + MEM[10637];
assign MEM[24727] = MEM[9430] + MEM[12543];
assign MEM[24728] = MEM[9438] + MEM[13309];
assign MEM[24729] = MEM[9440] + MEM[12128];
assign MEM[24730] = MEM[9442] + MEM[9650];
assign MEM[24731] = MEM[9444] + MEM[13045];
assign MEM[24732] = MEM[9450] + MEM[12458];
assign MEM[24733] = MEM[9453] + MEM[9536];
assign MEM[24734] = MEM[9466] + MEM[11792];
assign MEM[24735] = MEM[9468] + MEM[13291];
assign MEM[24736] = MEM[9473] + MEM[10811];
assign MEM[24737] = MEM[9476] + MEM[10403];
assign MEM[24738] = MEM[9479] + MEM[10046];
assign MEM[24739] = MEM[9486] + MEM[10175];
assign MEM[24740] = MEM[9488] + MEM[11614];
assign MEM[24741] = MEM[9495] + MEM[12568];
assign MEM[24742] = MEM[9501] + MEM[11885];
assign MEM[24743] = MEM[9506] + MEM[11136];
assign MEM[24744] = MEM[9507] + MEM[12662];
assign MEM[24745] = MEM[9518] + MEM[11940];
assign MEM[24746] = MEM[9522] + MEM[10368];
assign MEM[24747] = MEM[9525] + MEM[12596];
assign MEM[24748] = MEM[9530] + MEM[10732];
assign MEM[24749] = MEM[9535] + MEM[10306];
assign MEM[24750] = MEM[9544] + MEM[11509];
assign MEM[24751] = MEM[9551] + MEM[11796];
assign MEM[24752] = MEM[9555] + MEM[10696];
assign MEM[24753] = MEM[9563] + MEM[9869];
assign MEM[24754] = MEM[9568] + MEM[10147];
assign MEM[24755] = MEM[9582] + MEM[9992];
assign MEM[24756] = MEM[9587] + MEM[10426];
assign MEM[24757] = MEM[9588] + MEM[11121];
assign MEM[24758] = MEM[9610] + MEM[12430];
assign MEM[24759] = MEM[9615] + MEM[12285];
assign MEM[24760] = MEM[9616] + MEM[12449];
assign MEM[24761] = MEM[9617] + MEM[10506];
assign MEM[24762] = MEM[9617] + MEM[10955];
assign MEM[24763] = MEM[9628] + MEM[12001];
assign MEM[24764] = MEM[9636] + MEM[13921];
assign MEM[24765] = MEM[9637] + MEM[12435];
assign MEM[24766] = MEM[9646] + MEM[12561];
assign MEM[24767] = MEM[9648] + MEM[12107];
assign MEM[24768] = MEM[9653] + MEM[10264];
assign MEM[24769] = MEM[9675] + MEM[9809];
assign MEM[24770] = MEM[9683] + MEM[13775];
assign MEM[24771] = MEM[9709] + MEM[10785];
assign MEM[24772] = MEM[9717] + MEM[11318];
assign MEM[24773] = MEM[9735] + MEM[10221];
assign MEM[24774] = MEM[9739] + MEM[11795];
assign MEM[24775] = MEM[9747] + MEM[11581];
assign MEM[24776] = MEM[9750] + MEM[12215];
assign MEM[24777] = MEM[9770] + MEM[10024];
assign MEM[24778] = MEM[9773] + MEM[15270];
assign MEM[24779] = MEM[9796] + MEM[11892];
assign MEM[24780] = MEM[9805] + MEM[11567];
assign MEM[24781] = MEM[9840] + MEM[12142];
assign MEM[24782] = MEM[9841] + MEM[12454];
assign MEM[24783] = MEM[9862] + MEM[13640];
assign MEM[24784] = MEM[9870] + MEM[11539];
assign MEM[24785] = MEM[9880] + MEM[11763];
assign MEM[24786] = MEM[9888] + MEM[15498];
assign MEM[24787] = MEM[9890] + MEM[10945];
assign MEM[24788] = MEM[9898] + MEM[10593];
assign MEM[24789] = MEM[9900] + MEM[11901];
assign MEM[24790] = MEM[9901] + MEM[15201];
assign MEM[24791] = MEM[9905] + MEM[10586];
assign MEM[24792] = MEM[9916] + MEM[11046];
assign MEM[24793] = MEM[9942] + MEM[9985];
assign MEM[24794] = MEM[9948] + MEM[10062];
assign MEM[24795] = MEM[9953] + MEM[13672];
assign MEM[24796] = MEM[9957] + MEM[10337];
assign MEM[24797] = MEM[9968] + MEM[12246];
assign MEM[24798] = MEM[9970] + MEM[13083];
assign MEM[24799] = MEM[9976] + MEM[10054];
assign MEM[24800] = MEM[9981] + MEM[13072];
assign MEM[24801] = MEM[9988] + MEM[10780];
assign MEM[24802] = MEM[9994] + MEM[11977];
assign MEM[24803] = MEM[9998] + MEM[11152];
assign MEM[24804] = MEM[10001] + MEM[11556];
assign MEM[24805] = MEM[10033] + MEM[11834];
assign MEM[24806] = MEM[10038] + MEM[12117];
assign MEM[24807] = MEM[10040] + MEM[10665];
assign MEM[24808] = MEM[10059] + MEM[14152];
assign MEM[24809] = MEM[10062] + MEM[11595];
assign MEM[24810] = MEM[10083] + MEM[15975];
assign MEM[24811] = MEM[10084] + MEM[11710];
assign MEM[24812] = MEM[10098] + MEM[13667];
assign MEM[24813] = MEM[10109] + MEM[12151];
assign MEM[24814] = MEM[10111] + MEM[12773];
assign MEM[24815] = MEM[10112] + MEM[11465];
assign MEM[24816] = MEM[10114] + MEM[10206];
assign MEM[24817] = MEM[10119] + MEM[10886];
assign MEM[24818] = MEM[10122] + MEM[10392];
assign MEM[24819] = MEM[10125] + MEM[13769];
assign MEM[24820] = MEM[10128] + MEM[11766];
assign MEM[24821] = MEM[10130] + MEM[11149];
assign MEM[24822] = MEM[10134] + MEM[15689];
assign MEM[24823] = MEM[10143] + MEM[11478];
assign MEM[24824] = MEM[10145] + MEM[10149];
assign MEM[24825] = MEM[10151] + MEM[13335];
assign MEM[24826] = MEM[10156] + MEM[14346];
assign MEM[24827] = MEM[10163] + MEM[12119];
assign MEM[24828] = MEM[10173] + MEM[13150];
assign MEM[24829] = MEM[10179] + MEM[12346];
assign MEM[24830] = MEM[10182] + MEM[13655];
assign MEM[24831] = MEM[10190] + MEM[10910];
assign MEM[24832] = MEM[10194] + MEM[11845];
assign MEM[24833] = MEM[10197] + MEM[14812];
assign MEM[24834] = MEM[10208] + MEM[11658];
assign MEM[24835] = MEM[10217] + MEM[12149];
assign MEM[24836] = MEM[10218] + MEM[12130];
assign MEM[24837] = MEM[10220] + MEM[14260];
assign MEM[24838] = MEM[10245] + MEM[12344];
assign MEM[24839] = MEM[10247] + MEM[11701];
assign MEM[24840] = MEM[10248] + MEM[10901];
assign MEM[24841] = MEM[10248] + MEM[11685];
assign MEM[24842] = MEM[10250] + MEM[14572];
assign MEM[24843] = MEM[10257] + MEM[11056];
assign MEM[24844] = MEM[10260] + MEM[10826];
assign MEM[24845] = MEM[10275] + MEM[10710];
assign MEM[24846] = MEM[10286] + MEM[12618];
assign MEM[24847] = MEM[10288] + MEM[11839];
assign MEM[24848] = MEM[10304] + MEM[10532];
assign MEM[24849] = MEM[10307] + MEM[10783];
assign MEM[24850] = MEM[10309] + MEM[13552];
assign MEM[24851] = MEM[10318] + MEM[10523];
assign MEM[24852] = MEM[10320] + MEM[11093];
assign MEM[24853] = MEM[10330] + MEM[13230];
assign MEM[24854] = MEM[10332] + MEM[11950];
assign MEM[24855] = MEM[10333] + MEM[11139];
assign MEM[24856] = MEM[10345] + MEM[10755];
assign MEM[24857] = MEM[10350] + MEM[10448];
assign MEM[24858] = MEM[10351] + MEM[11610];
assign MEM[24859] = MEM[10354] + MEM[12630];
assign MEM[24860] = MEM[10373] + MEM[12762];
assign MEM[24861] = MEM[10382] + MEM[11990];
assign MEM[24862] = MEM[10383] + MEM[12267];
assign MEM[24863] = MEM[10391] + MEM[10711];
assign MEM[24864] = MEM[10405] + MEM[10761];
assign MEM[24865] = MEM[10415] + MEM[10928];
assign MEM[24866] = MEM[10417] + MEM[12700];
assign MEM[24867] = MEM[10427] + MEM[13483];
assign MEM[24868] = MEM[10431] + MEM[11004];
assign MEM[24869] = MEM[10435] + MEM[10498];
assign MEM[24870] = MEM[10435] + MEM[15417];
assign MEM[24871] = MEM[10439] + MEM[12384];
assign MEM[24872] = MEM[10444] + MEM[13300];
assign MEM[24873] = MEM[10459] + MEM[15442];
assign MEM[24874] = MEM[10460] + MEM[10522];
assign MEM[24875] = MEM[10463] + MEM[12099];
assign MEM[24876] = MEM[10474] + MEM[12520];
assign MEM[24877] = MEM[10475] + MEM[16007];
assign MEM[24878] = MEM[10479] + MEM[11544];
assign MEM[24879] = MEM[10480] + MEM[11010];
assign MEM[24880] = MEM[10483] + MEM[11572];
assign MEM[24881] = MEM[10503] + MEM[14104];
assign MEM[24882] = MEM[10515] + MEM[12575];
assign MEM[24883] = MEM[10518] + MEM[11922];
assign MEM[24884] = MEM[10520] + MEM[10748];
assign MEM[24885] = MEM[10526] + MEM[11916];
assign MEM[24886] = MEM[10527] + MEM[11628];
assign MEM[24887] = MEM[10535] + MEM[11677];
assign MEM[24888] = MEM[10551] + MEM[11693];
assign MEM[24889] = MEM[10554] + MEM[12659];
assign MEM[24890] = MEM[10555] + MEM[13006];
assign MEM[24891] = MEM[10566] + MEM[11035];
assign MEM[24892] = MEM[10571] + MEM[13002];
assign MEM[24893] = MEM[10572] + MEM[11213];
assign MEM[24894] = MEM[10573] + MEM[10676];
assign MEM[24895] = MEM[10583] + MEM[11006];
assign MEM[24896] = MEM[10587] + MEM[11625];
assign MEM[24897] = MEM[10592] + MEM[12173];
assign MEM[24898] = MEM[10599] + MEM[14456];
assign MEM[24899] = MEM[10605] + MEM[10740];
assign MEM[24900] = MEM[10610] + MEM[11919];
assign MEM[24901] = MEM[10613] + MEM[13047];
assign MEM[24902] = MEM[10614] + MEM[12730];
assign MEM[24903] = MEM[10622] + MEM[11537];
assign MEM[24904] = MEM[10626] + MEM[11936];
assign MEM[24905] = MEM[10628] + MEM[16484];
assign MEM[24906] = MEM[10630] + MEM[17816];
assign MEM[24907] = MEM[10632] + MEM[11615];
assign MEM[24908] = MEM[10635] + MEM[12064];
assign MEM[24909] = MEM[10638] + MEM[10771];
assign MEM[24910] = MEM[10641] + MEM[14793];
assign MEM[24911] = MEM[10642] + MEM[12437];
assign MEM[24912] = MEM[10646] + MEM[10878];
assign MEM[24913] = MEM[10650] + MEM[10987];
assign MEM[24914] = MEM[10651] + MEM[15089];
assign MEM[24915] = MEM[10652] + MEM[13348];
assign MEM[24916] = MEM[10653] + MEM[15080];
assign MEM[24917] = MEM[10655] + MEM[10674];
assign MEM[24918] = MEM[10657] + MEM[13350];
assign MEM[24919] = MEM[10660] + MEM[13263];
assign MEM[24920] = MEM[10662] + MEM[11249];
assign MEM[24921] = MEM[10669] + MEM[11897];
assign MEM[24922] = MEM[10679] + MEM[12827];
assign MEM[24923] = MEM[10680] + MEM[12171];
assign MEM[24924] = MEM[10681] + MEM[11031];
assign MEM[24925] = MEM[10688] + MEM[15424];
assign MEM[24926] = MEM[10698] + MEM[15512];
assign MEM[24927] = MEM[10700] + MEM[11653];
assign MEM[24928] = MEM[10701] + MEM[14656];
assign MEM[24929] = MEM[10704] + MEM[11203];
assign MEM[24930] = MEM[10706] + MEM[10973];
assign MEM[24931] = MEM[10707] + MEM[13500];
assign MEM[24932] = MEM[10709] + MEM[12869];
assign MEM[24933] = MEM[10713] + MEM[13965];
assign MEM[24934] = MEM[10714] + MEM[14659];
assign MEM[24935] = MEM[10715] + MEM[11126];
assign MEM[24936] = MEM[10719] + MEM[13419];
assign MEM[24937] = MEM[10724] + MEM[11985];
assign MEM[24938] = MEM[10727] + MEM[12410];
assign MEM[24939] = MEM[10729] + MEM[11832];
assign MEM[24940] = MEM[10730] + MEM[11266];
assign MEM[24941] = MEM[10731] + MEM[11184];
assign MEM[24942] = MEM[10737] + MEM[11312];
assign MEM[24943] = MEM[10738] + MEM[13212];
assign MEM[24944] = MEM[10744] + MEM[16762];
assign MEM[24945] = MEM[10745] + MEM[12868];
assign MEM[24946] = MEM[10753] + MEM[13068];
assign MEM[24947] = MEM[10756] + MEM[10976];
assign MEM[24948] = MEM[10765] + MEM[10882];
assign MEM[24949] = MEM[10766] + MEM[12145];
assign MEM[24950] = MEM[10768] + MEM[13165];
assign MEM[24951] = MEM[10769] + MEM[14546];
assign MEM[24952] = MEM[10773] + MEM[10846];
assign MEM[24953] = MEM[10777] + MEM[12538];
assign MEM[24954] = MEM[10778] + MEM[11793];
assign MEM[24955] = MEM[10781] + MEM[13204];
assign MEM[24956] = MEM[10784] + MEM[19755];
assign MEM[24957] = MEM[10788] + MEM[12369];
assign MEM[24958] = MEM[10788] + MEM[13574];
assign MEM[24959] = MEM[10789] + MEM[11679];
assign MEM[24960] = MEM[10792] + MEM[10929];
assign MEM[24961] = MEM[10793] + MEM[12979];
assign MEM[24962] = MEM[10795] + MEM[12353];
assign MEM[24963] = MEM[10796] + MEM[11995];
assign MEM[24964] = MEM[10797] + MEM[11838];
assign MEM[24965] = MEM[10798] + MEM[13457];
assign MEM[24966] = MEM[10799] + MEM[12930];
assign MEM[24967] = MEM[10807] + MEM[12154];
assign MEM[24968] = MEM[10808] + MEM[13255];
assign MEM[24969] = MEM[10809] + MEM[11690];
assign MEM[24970] = MEM[10810] + MEM[13825];
assign MEM[24971] = MEM[10812] + MEM[12746];
assign MEM[24972] = MEM[10819] + MEM[12935];
assign MEM[24973] = MEM[10820] + MEM[12150];
assign MEM[24974] = MEM[10821] + MEM[14080];
assign MEM[24975] = MEM[10824] + MEM[12238];
assign MEM[24976] = MEM[10825] + MEM[13602];
assign MEM[24977] = MEM[10829] + MEM[11787];
assign MEM[24978] = MEM[10830] + MEM[11890];
assign MEM[24979] = MEM[10832] + MEM[13523];
assign MEM[24980] = MEM[10834] + MEM[12617];
assign MEM[24981] = MEM[10835] + MEM[13848];
assign MEM[24982] = MEM[10837] + MEM[12376];
assign MEM[24983] = MEM[10838] + MEM[16516];
assign MEM[24984] = MEM[10840] + MEM[10978];
assign MEM[24985] = MEM[10843] + MEM[11464];
assign MEM[24986] = MEM[10848] + MEM[15999];
assign MEM[24987] = MEM[10849] + MEM[12260];
assign MEM[24988] = MEM[10850] + MEM[12977];
assign MEM[24989] = MEM[10851] + MEM[12125];
assign MEM[24990] = MEM[10854] + MEM[12505];
assign MEM[24991] = MEM[10857] + MEM[13282];
assign MEM[24992] = MEM[10858] + MEM[11826];
assign MEM[24993] = MEM[10867] + MEM[11599];
assign MEM[24994] = MEM[10871] + MEM[11172];
assign MEM[24995] = MEM[10872] + MEM[12081];
assign MEM[24996] = MEM[10874] + MEM[12534];
assign MEM[24997] = MEM[10877] + MEM[15265];
assign MEM[24998] = MEM[10879] + MEM[13422];
assign MEM[24999] = MEM[10881] + MEM[12620];
assign MEM[25000] = MEM[10883] + MEM[12061];
assign MEM[25001] = MEM[10885] + MEM[13897];
assign MEM[25002] = MEM[10893] + MEM[14800];
assign MEM[25003] = MEM[10897] + MEM[12582];
assign MEM[25004] = MEM[10898] + MEM[12301];
assign MEM[25005] = MEM[10899] + MEM[10903];
assign MEM[25006] = MEM[10900] + MEM[11530];
assign MEM[25007] = MEM[10904] + MEM[12153];
assign MEM[25008] = MEM[10905] + MEM[14540];
assign MEM[25009] = MEM[10906] + MEM[12336];
assign MEM[25010] = MEM[10911] + MEM[11700];
assign MEM[25011] = MEM[10916] + MEM[11028];
assign MEM[25012] = MEM[10919] + MEM[13017];
assign MEM[25013] = MEM[10920] + MEM[11837];
assign MEM[25014] = MEM[10921] + MEM[12510];
assign MEM[25015] = MEM[10922] + MEM[14854];
assign MEM[25016] = MEM[10925] + MEM[15939];
assign MEM[25017] = MEM[10926] + MEM[10934];
assign MEM[25018] = MEM[10930] + MEM[11304];
assign MEM[25019] = MEM[10935] + MEM[12950];
assign MEM[25020] = MEM[10939] + MEM[13184];
assign MEM[25021] = MEM[10940] + MEM[12293];
assign MEM[25022] = MEM[10946] + MEM[11652];
assign MEM[25023] = MEM[10947] + MEM[12855];
assign MEM[25024] = MEM[10948] + MEM[13351];
assign MEM[25025] = MEM[10950] + MEM[12484];
assign MEM[25026] = MEM[10956] + MEM[12091];
assign MEM[25027] = MEM[10958] + MEM[11775];
assign MEM[25028] = MEM[10961] + MEM[16536];
assign MEM[25029] = MEM[10963] + MEM[12187];
assign MEM[25030] = MEM[10966] + MEM[11666];
assign MEM[25031] = MEM[10968] + MEM[13182];
assign MEM[25032] = MEM[10970] + MEM[11022];
assign MEM[25033] = MEM[10972] + MEM[11106];
assign MEM[25034] = MEM[10974] + MEM[11110];
assign MEM[25035] = MEM[10975] + MEM[12002];
assign MEM[25036] = MEM[10977] + MEM[11632];
assign MEM[25037] = MEM[10979] + MEM[15845];
assign MEM[25038] = MEM[10980] + MEM[14705];
assign MEM[25039] = MEM[10981] + MEM[12968];
assign MEM[25040] = MEM[10985] + MEM[16066];
assign MEM[25041] = MEM[10986] + MEM[13244];
assign MEM[25042] = MEM[10988] + MEM[11027];
assign MEM[25043] = MEM[10992] + MEM[11780];
assign MEM[25044] = MEM[10993] + MEM[14755];
assign MEM[25045] = MEM[10996] + MEM[12556];
assign MEM[25046] = MEM[10997] + MEM[14210];
assign MEM[25047] = MEM[11003] + MEM[11406];
assign MEM[25048] = MEM[11005] + MEM[11101];
assign MEM[25049] = MEM[11012] + MEM[11016];
assign MEM[25050] = MEM[11023] + MEM[13474];
assign MEM[25051] = MEM[11026] + MEM[15520];
assign MEM[25052] = MEM[11030] + MEM[13012];
assign MEM[25053] = MEM[11032] + MEM[13968];
assign MEM[25054] = MEM[11037] + MEM[11755];
assign MEM[25055] = MEM[11040] + MEM[12462];
assign MEM[25056] = MEM[11041] + MEM[12976];
assign MEM[25057] = MEM[11042] + MEM[14587];
assign MEM[25058] = MEM[11048] + MEM[14175];
assign MEM[25059] = MEM[11052] + MEM[12020];
assign MEM[25060] = MEM[11054] + MEM[13594];
assign MEM[25061] = MEM[11055] + MEM[12720];
assign MEM[25062] = MEM[11057] + MEM[11745];
assign MEM[25063] = MEM[11059] + MEM[12405];
assign MEM[25064] = MEM[11060] + MEM[15051];
assign MEM[25065] = MEM[11061] + MEM[11255];
assign MEM[25066] = MEM[11062] + MEM[11992];
assign MEM[25067] = MEM[11063] + MEM[12969];
assign MEM[25068] = MEM[11064] + MEM[12122];
assign MEM[25069] = MEM[11065] + MEM[11083];
assign MEM[25070] = MEM[11069] + MEM[16247];
assign MEM[25071] = MEM[11072] + MEM[12711];
assign MEM[25072] = MEM[11075] + MEM[12050];
assign MEM[25073] = MEM[11077] + MEM[11866];
assign MEM[25074] = MEM[11078] + MEM[12186];
assign MEM[25075] = MEM[11079] + MEM[12625];
assign MEM[25076] = MEM[11090] + MEM[12280];
assign MEM[25077] = MEM[11091] + MEM[12588];
assign MEM[25078] = MEM[11096] + MEM[11622];
assign MEM[25079] = MEM[11098] + MEM[12025];
assign MEM[25080] = MEM[11102] + MEM[15547];
assign MEM[25081] = MEM[11112] + MEM[16997];
assign MEM[25082] = MEM[11113] + MEM[16203];
assign MEM[25083] = MEM[11114] + MEM[11295];
assign MEM[25084] = MEM[11115] + MEM[12195];
assign MEM[25085] = MEM[11118] + MEM[16367];
assign MEM[25086] = MEM[11119] + MEM[17237];
assign MEM[25087] = MEM[11123] + MEM[12531];
assign MEM[25088] = MEM[11127] + MEM[14790];
assign MEM[25089] = MEM[11128] + MEM[13257];
assign MEM[25090] = MEM[11130] + MEM[15298];
assign MEM[25091] = MEM[11134] + MEM[15241];
assign MEM[25092] = MEM[11138] + MEM[11934];
assign MEM[25093] = MEM[11140] + MEM[11616];
assign MEM[25094] = MEM[11141] + MEM[14408];
assign MEM[25095] = MEM[11143] + MEM[11237];
assign MEM[25096] = MEM[11144] + MEM[13536];
assign MEM[25097] = MEM[11147] + MEM[14207];
assign MEM[25098] = MEM[11148] + MEM[11967];
assign MEM[25099] = MEM[11150] + MEM[11326];
assign MEM[25100] = MEM[11153] + MEM[13929];
assign MEM[25101] = MEM[11154] + MEM[12427];
assign MEM[25102] = MEM[11158] + MEM[16434];
assign MEM[25103] = MEM[11159] + MEM[12180];
assign MEM[25104] = MEM[11160] + MEM[15332];
assign MEM[25105] = MEM[11161] + MEM[11854];
assign MEM[25106] = MEM[11163] + MEM[12439];
assign MEM[25107] = MEM[11164] + MEM[12587];
assign MEM[25108] = MEM[11167] + MEM[14366];
assign MEM[25109] = MEM[11171] + MEM[13228];
assign MEM[25110] = MEM[11177] + MEM[12581];
assign MEM[25111] = MEM[11178] + MEM[12432];
assign MEM[25112] = MEM[11179] + MEM[13429];
assign MEM[25113] = MEM[11181] + MEM[13079];
assign MEM[25114] = MEM[11183] + MEM[12343];
assign MEM[25115] = MEM[11185] + MEM[13283];
assign MEM[25116] = MEM[11186] + MEM[11806];
assign MEM[25117] = MEM[11190] + MEM[12877];
assign MEM[25118] = MEM[11193] + MEM[15327];
assign MEM[25119] = MEM[11195] + MEM[14916];
assign MEM[25120] = MEM[11210] + MEM[11212];
assign MEM[25121] = MEM[11212] + MEM[13007];
assign MEM[25122] = MEM[11214] + MEM[15096];
assign MEM[25123] = MEM[11215] + MEM[14894];
assign MEM[25124] = MEM[11217] + MEM[12497];
assign MEM[25125] = MEM[11218] + MEM[14584];
assign MEM[25126] = MEM[11219] + MEM[12854];
assign MEM[25127] = MEM[11222] + MEM[11274];
assign MEM[25128] = MEM[11223] + MEM[11328];
assign MEM[25129] = MEM[11226] + MEM[14208];
assign MEM[25130] = MEM[11228] + MEM[13557];
assign MEM[25131] = MEM[11229] + MEM[13829];
assign MEM[25132] = MEM[11231] + MEM[11833];
assign MEM[25133] = MEM[11233] + MEM[11502];
assign MEM[25134] = MEM[11238] + MEM[14453];
assign MEM[25135] = MEM[11248] + MEM[11864];
assign MEM[25136] = MEM[11254] + MEM[11596];
assign MEM[25137] = MEM[11256] + MEM[14205];
assign MEM[25138] = MEM[11258] + MEM[12571];
assign MEM[25139] = MEM[11265] + MEM[16342];
assign MEM[25140] = MEM[11276] + MEM[15578];
assign MEM[25141] = MEM[11278] + MEM[19771];
assign MEM[25142] = MEM[11280] + MEM[15439];
assign MEM[25143] = MEM[11282] + MEM[11751];
assign MEM[25144] = MEM[11284] + MEM[13580];
assign MEM[25145] = MEM[11291] + MEM[12631];
assign MEM[25146] = MEM[11292] + MEM[13042];
assign MEM[25147] = MEM[11293] + MEM[12057];
assign MEM[25148] = MEM[11294] + MEM[12816];
assign MEM[25149] = MEM[11299] + MEM[13666];
assign MEM[25150] = MEM[11300] + MEM[11960];
assign MEM[25151] = MEM[11307] + MEM[12738];
assign MEM[25152] = MEM[11308] + MEM[13865];
assign MEM[25153] = MEM[11320] + MEM[12989];
assign MEM[25154] = MEM[11323] + MEM[14797];
assign MEM[25155] = MEM[11327] + MEM[16867];
assign MEM[25156] = MEM[11345] + MEM[13372];
assign MEM[25157] = MEM[11354] + MEM[11640];
assign MEM[25158] = MEM[11357] + MEM[11583];
assign MEM[25159] = MEM[11375] + MEM[13780];
assign MEM[25160] = MEM[11381] + MEM[11554];
assign MEM[25161] = MEM[11391] + MEM[12075];
assign MEM[25162] = MEM[11406] + MEM[16521];
assign MEM[25163] = MEM[11422] + MEM[12842];
assign MEM[25164] = MEM[11431] + MEM[11844];
assign MEM[25165] = MEM[11443] + MEM[12136];
assign MEM[25166] = MEM[11456] + MEM[11743];
assign MEM[25167] = MEM[11459] + MEM[11933];
assign MEM[25168] = MEM[11483] + MEM[13533];
assign MEM[25169] = MEM[11501] + MEM[14044];
assign MEM[25170] = MEM[11543] + MEM[12886];
assign MEM[25171] = MEM[11550] + MEM[13019];
assign MEM[25172] = MEM[11565] + MEM[11735];
assign MEM[25173] = MEM[11573] + MEM[12089];
assign MEM[25174] = MEM[11589] + MEM[14112];
assign MEM[25175] = MEM[11602] + MEM[12431];
assign MEM[25176] = MEM[11605] + MEM[12882];
assign MEM[25177] = MEM[11608] + MEM[11784];
assign MEM[25178] = MEM[11609] + MEM[13637];
assign MEM[25179] = MEM[11613] + MEM[12453];
assign MEM[25180] = MEM[11621] + MEM[12761];
assign MEM[25181] = MEM[11624] + MEM[12313];
assign MEM[25182] = MEM[11638] + MEM[12361];
assign MEM[25183] = MEM[11639] + MEM[13280];
assign MEM[25184] = MEM[11665] + MEM[12515];
assign MEM[25185] = MEM[11669] + MEM[11848];
assign MEM[25186] = MEM[11675] + MEM[12059];
assign MEM[25187] = MEM[11707] + MEM[13634];
assign MEM[25188] = MEM[11714] + MEM[11893];
assign MEM[25189] = MEM[11714] + MEM[12468];
assign MEM[25190] = MEM[11725] + MEM[12212];
assign MEM[25191] = MEM[11730] + MEM[12553];
assign MEM[25192] = MEM[11737] + MEM[11898];
assign MEM[25193] = MEM[11741] + MEM[11876];
assign MEM[25194] = MEM[11744] + MEM[12595];
assign MEM[25195] = MEM[11752] + MEM[12192];
assign MEM[25196] = MEM[11782] + MEM[12067];
assign MEM[25197] = MEM[11790] + MEM[13383];
assign MEM[25198] = MEM[11798] + MEM[12417];
assign MEM[25199] = MEM[11813] + MEM[12068];
assign MEM[25200] = MEM[11817] + MEM[11942];
assign MEM[25201] = MEM[11819] + MEM[12236];
assign MEM[25202] = MEM[11841] + MEM[12765];
assign MEM[25203] = MEM[11849] + MEM[13349];
assign MEM[25204] = MEM[11862] + MEM[12191];
assign MEM[25205] = MEM[11865] + MEM[12110];
assign MEM[25206] = MEM[11867] + MEM[12440];
assign MEM[25207] = MEM[11873] + MEM[14610];
assign MEM[25208] = MEM[11883] + MEM[12209];
assign MEM[25209] = MEM[11887] + MEM[12258];
assign MEM[25210] = MEM[11889] + MEM[13107];
assign MEM[25211] = MEM[11905] + MEM[12768];
assign MEM[25212] = MEM[11907] + MEM[12314];
assign MEM[25213] = MEM[11910] + MEM[15253];
assign MEM[25214] = MEM[11914] + MEM[12086];
assign MEM[25215] = MEM[11931] + MEM[12902];
assign MEM[25216] = MEM[11932] + MEM[12812];
assign MEM[25217] = MEM[11935] + MEM[13440];
assign MEM[25218] = MEM[11937] + MEM[12374];
assign MEM[25219] = MEM[11938] + MEM[13932];
assign MEM[25220] = MEM[11944] + MEM[12729];
assign MEM[25221] = MEM[11945] + MEM[13541];
assign MEM[25222] = MEM[11946] + MEM[12098];
assign MEM[25223] = MEM[11957] + MEM[12201];
assign MEM[25224] = MEM[11958] + MEM[12574];
assign MEM[25225] = MEM[11959] + MEM[12302];
assign MEM[25226] = MEM[11965] + MEM[13678];
assign MEM[25227] = MEM[11969] + MEM[12887];
assign MEM[25228] = MEM[11982] + MEM[12477];
assign MEM[25229] = MEM[11989] + MEM[12311];
assign MEM[25230] = MEM[11993] + MEM[12604];
assign MEM[25231] = MEM[11997] + MEM[12170];
assign MEM[25232] = MEM[11998] + MEM[12638];
assign MEM[25233] = MEM[11998] + MEM[14074];
assign MEM[25234] = MEM[12009] + MEM[12271];
assign MEM[25235] = MEM[12011] + MEM[13271];
assign MEM[25236] = MEM[12019] + MEM[12493];
assign MEM[25237] = MEM[12020] + MEM[12988];
assign MEM[25238] = MEM[12037] + MEM[12452];
assign MEM[25239] = MEM[12047] + MEM[12649];
assign MEM[25240] = MEM[12058] + MEM[14075];
assign MEM[25241] = MEM[12060] + MEM[12211];
assign MEM[25242] = MEM[12067] + MEM[16021];
assign MEM[25243] = MEM[12070] + MEM[12159];
assign MEM[25244] = MEM[12073] + MEM[12438];
assign MEM[25245] = MEM[12074] + MEM[14514];
assign MEM[25246] = MEM[12085] + MEM[14017];
assign MEM[25247] = MEM[12087] + MEM[12564];
assign MEM[25248] = MEM[12090] + MEM[12179];
assign MEM[25249] = MEM[12093] + MEM[13363];
assign MEM[25250] = MEM[12094] + MEM[15893];
assign MEM[25251] = MEM[12095] + MEM[13090];
assign MEM[25252] = MEM[12096] + MEM[16389];
assign MEM[25253] = MEM[12097] + MEM[15910];
assign MEM[25254] = MEM[12101] + MEM[12210];
assign MEM[25255] = MEM[12104] + MEM[12295];
assign MEM[25256] = MEM[12105] + MEM[13270];
assign MEM[25257] = MEM[12111] + MEM[16085];
assign MEM[25258] = MEM[12112] + MEM[14144];
assign MEM[25259] = MEM[12114] + MEM[12763];
assign MEM[25260] = MEM[12115] + MEM[13441];
assign MEM[25261] = MEM[12120] + MEM[15230];
assign MEM[25262] = MEM[12123] + MEM[16650];
assign MEM[25263] = MEM[12124] + MEM[15625];
assign MEM[25264] = MEM[12127] + MEM[12962];
assign MEM[25265] = MEM[12129] + MEM[12905];
assign MEM[25266] = MEM[12131] + MEM[17284];
assign MEM[25267] = MEM[12132] + MEM[14937];
assign MEM[25268] = MEM[12134] + MEM[12402];
assign MEM[25269] = MEM[12135] + MEM[12200];
assign MEM[25270] = MEM[12140] + MEM[12365];
assign MEM[25271] = MEM[12141] + MEM[13113];
assign MEM[25272] = MEM[12143] + MEM[12483];
assign MEM[25273] = MEM[12155] + MEM[13367];
assign MEM[25274] = MEM[12158] + MEM[13293];
assign MEM[25275] = MEM[12160] + MEM[12290];
assign MEM[25276] = MEM[12164] + MEM[12373];
assign MEM[25277] = MEM[12167] + MEM[13317];
assign MEM[25278] = MEM[12168] + MEM[12172];
assign MEM[25279] = MEM[12169] + MEM[14685];
assign MEM[25280] = MEM[12175] + MEM[13463];
assign MEM[25281] = MEM[12176] + MEM[14385];
assign MEM[25282] = MEM[12177] + MEM[13700];
assign MEM[25283] = MEM[12178] + MEM[16293];
assign MEM[25284] = MEM[12181] + MEM[16914];
assign MEM[25285] = MEM[12190] + MEM[13357];
assign MEM[25286] = MEM[12193] + MEM[17401];
assign MEM[25287] = MEM[12194] + MEM[12642];
assign MEM[25288] = MEM[12197] + MEM[14095];
assign MEM[25289] = MEM[12198] + MEM[18592];
assign MEM[25290] = MEM[12202] + MEM[12602];
assign MEM[25291] = MEM[12203] + MEM[12521];
assign MEM[25292] = MEM[12204] + MEM[18119];
assign MEM[25293] = MEM[12207] + MEM[13779];
assign MEM[25294] = MEM[12208] + MEM[12972];
assign MEM[25295] = MEM[12213] + MEM[12743];
assign MEM[25296] = MEM[12214] + MEM[15299];
assign MEM[25297] = MEM[12217] + MEM[16190];
assign MEM[25298] = MEM[12221] + MEM[12433];
assign MEM[25299] = MEM[12223] + MEM[13787];
assign MEM[25300] = MEM[12224] + MEM[13890];
assign MEM[25301] = MEM[12226] + MEM[13418];
assign MEM[25302] = MEM[12229] + MEM[15041];
assign MEM[25303] = MEM[12230] + MEM[13799];
assign MEM[25304] = MEM[12233] + MEM[16509];
assign MEM[25305] = MEM[12234] + MEM[12249];
assign MEM[25306] = MEM[12237] + MEM[12456];
assign MEM[25307] = MEM[12241] + MEM[12707];
assign MEM[25308] = MEM[12243] + MEM[15627];
assign MEM[25309] = MEM[12251] + MEM[14295];
assign MEM[25310] = MEM[12253] + MEM[12600];
assign MEM[25311] = MEM[12254] + MEM[13938];
assign MEM[25312] = MEM[12255] + MEM[13777];
assign MEM[25313] = MEM[12257] + MEM[12611];
assign MEM[25314] = MEM[12262] + MEM[13246];
assign MEM[25315] = MEM[12264] + MEM[14096];
assign MEM[25316] = MEM[12266] + MEM[14221];
assign MEM[25317] = MEM[12270] + MEM[13149];
assign MEM[25318] = MEM[12274] + MEM[17058];
assign MEM[25319] = MEM[12275] + MEM[15937];
assign MEM[25320] = MEM[12279] + MEM[13527];
assign MEM[25321] = MEM[12287] + MEM[12705];
assign MEM[25322] = MEM[12289] + MEM[13583];
assign MEM[25323] = MEM[12291] + MEM[17185];
assign MEM[25324] = MEM[12304] + MEM[13420];
assign MEM[25325] = MEM[12305] + MEM[15790];
assign MEM[25326] = MEM[12306] + MEM[12819];
assign MEM[25327] = MEM[12307] + MEM[17190];
assign MEM[25328] = MEM[12310] + MEM[12970];
assign MEM[25329] = MEM[12315] + MEM[15206];
assign MEM[25330] = MEM[12316] + MEM[15750];
assign MEM[25331] = MEM[12317] + MEM[13569];
assign MEM[25332] = MEM[12320] + MEM[13426];
assign MEM[25333] = MEM[12323] + MEM[14970];
assign MEM[25334] = MEM[12326] + MEM[17180];
assign MEM[25335] = MEM[12328] + MEM[12948];
assign MEM[25336] = MEM[12330] + MEM[15666];
assign MEM[25337] = MEM[12332] + MEM[13919];
assign MEM[25338] = MEM[12338] + MEM[13702];
assign MEM[25339] = MEM[12339] + MEM[14428];
assign MEM[25340] = MEM[12348] + MEM[13140];
assign MEM[25341] = MEM[12352] + MEM[13392];
assign MEM[25342] = MEM[12354] + MEM[13381];
assign MEM[25343] = MEM[12355] + MEM[13234];
assign MEM[25344] = MEM[12357] + MEM[13338];
assign MEM[25345] = MEM[12358] + MEM[12863];
assign MEM[25346] = MEM[12371] + MEM[12379];
assign MEM[25347] = MEM[12372] + MEM[14342];
assign MEM[25348] = MEM[12377] + MEM[14227];
assign MEM[25349] = MEM[12378] + MEM[16363];
assign MEM[25350] = MEM[12382] + MEM[14933];
assign MEM[25351] = MEM[12383] + MEM[13688];
assign MEM[25352] = MEM[12385] + MEM[12416];
assign MEM[25353] = MEM[12390] + MEM[13156];
assign MEM[25354] = MEM[12392] + MEM[18174];
assign MEM[25355] = MEM[12396] + MEM[15760];
assign MEM[25356] = MEM[12398] + MEM[13129];
assign MEM[25357] = MEM[12399] + MEM[12668];
assign MEM[25358] = MEM[12403] + MEM[12678];
assign MEM[25359] = MEM[12404] + MEM[14444];
assign MEM[25360] = MEM[12406] + MEM[15049];
assign MEM[25361] = MEM[12409] + MEM[13509];
assign MEM[25362] = MEM[12411] + MEM[14601];
assign MEM[25363] = MEM[12412] + MEM[15923];
assign MEM[25364] = MEM[12415] + MEM[17498];
assign MEM[25365] = MEM[12419] + MEM[13209];
assign MEM[25366] = MEM[12420] + MEM[12963];
assign MEM[25367] = MEM[12421] + MEM[15417];
assign MEM[25368] = MEM[12422] + MEM[12526];
assign MEM[25369] = MEM[12423] + MEM[13375];
assign MEM[25370] = MEM[12428] + MEM[12633];
assign MEM[25371] = MEM[12429] + MEM[13088];
assign MEM[25372] = MEM[12434] + MEM[15624];
assign MEM[25373] = MEM[12436] + MEM[13241];
assign MEM[25374] = MEM[12441] + MEM[14409];
assign MEM[25375] = MEM[12442] + MEM[13644];
assign MEM[25376] = MEM[12443] + MEM[13674];
assign MEM[25377] = MEM[12445] + MEM[12805];
assign MEM[25378] = MEM[12451] + MEM[12971];
assign MEM[25379] = MEM[12457] + MEM[14417];
assign MEM[25380] = MEM[12459] + MEM[13412];
assign MEM[25381] = MEM[12461] + MEM[14167];
assign MEM[25382] = MEM[12464] + MEM[12921];
assign MEM[25383] = MEM[12466] + MEM[13195];
assign MEM[25384] = MEM[12467] + MEM[17170];
assign MEM[25385] = MEM[12470] + MEM[12793];
assign MEM[25386] = MEM[12471] + MEM[13373];
assign MEM[25387] = MEM[12475] + MEM[14080];
assign MEM[25388] = MEM[12479] + MEM[14284];
assign MEM[25389] = MEM[12481] + MEM[15793];
assign MEM[25390] = MEM[12486] + MEM[16117];
assign MEM[25391] = MEM[12488] + MEM[12641];
assign MEM[25392] = MEM[12489] + MEM[13835];
assign MEM[25393] = MEM[12490] + MEM[14604];
assign MEM[25394] = MEM[12491] + MEM[13022];
assign MEM[25395] = MEM[12492] + MEM[14515];
assign MEM[25396] = MEM[12496] + MEM[17279];
assign MEM[25397] = MEM[12502] + MEM[14379];
assign MEM[25398] = MEM[12503] + MEM[18510];
assign MEM[25399] = MEM[12507] + MEM[14741];
assign MEM[25400] = MEM[12508] + MEM[12551];
assign MEM[25401] = MEM[12511] + MEM[12590];
assign MEM[25402] = MEM[12513] + MEM[13461];
assign MEM[25403] = MEM[12516] + MEM[12589];
assign MEM[25404] = MEM[12517] + MEM[13397];
assign MEM[25405] = MEM[12519] + MEM[13223];
assign MEM[25406] = MEM[12522] + MEM[12903];
assign MEM[25407] = MEM[12523] + MEM[13478];
assign MEM[25408] = MEM[12527] + MEM[12766];
assign MEM[25409] = MEM[12529] + MEM[13442];
assign MEM[25410] = MEM[12530] + MEM[13809];
assign MEM[25411] = MEM[12532] + MEM[14238];
assign MEM[25412] = MEM[12539] + MEM[14069];
assign MEM[25413] = MEM[12540] + MEM[15635];
assign MEM[25414] = MEM[12542] + MEM[13824];
assign MEM[25415] = MEM[12545] + MEM[15489];
assign MEM[25416] = MEM[12546] + MEM[12567];
assign MEM[25417] = MEM[12547] + MEM[13370];
assign MEM[25418] = MEM[12548] + MEM[12736];
assign MEM[25419] = MEM[12549] + MEM[15861];
assign MEM[25420] = MEM[12552] + MEM[16702];
assign MEM[25421] = MEM[12554] + MEM[12821];
assign MEM[25422] = MEM[12559] + MEM[13652];
assign MEM[25423] = MEM[12563] + MEM[12628];
assign MEM[25424] = MEM[12569] + MEM[12978];
assign MEM[25425] = MEM[12570] + MEM[16400];
assign MEM[25426] = MEM[12572] + MEM[13104];
assign MEM[25427] = MEM[12579] + MEM[17934];
assign MEM[25428] = MEM[12585] + MEM[18669];
assign MEM[25429] = MEM[12592] + MEM[13029];
assign MEM[25430] = MEM[12597] + MEM[13119];
assign MEM[25431] = MEM[12598] + MEM[13589];
assign MEM[25432] = MEM[12601] + MEM[14363];
assign MEM[25433] = MEM[12603] + MEM[14785];
assign MEM[25434] = MEM[12605] + MEM[13559];
assign MEM[25435] = MEM[12606] + MEM[15771];
assign MEM[25436] = MEM[12607] + MEM[12704];
assign MEM[25437] = MEM[12608] + MEM[13122];
assign MEM[25438] = MEM[12609] + MEM[16388];
assign MEM[25439] = MEM[12613] + MEM[13028];
assign MEM[25440] = MEM[12614] + MEM[13586];
assign MEM[25441] = MEM[12615] + MEM[13287];
assign MEM[25442] = MEM[12616] + MEM[13054];
assign MEM[25443] = MEM[12621] + MEM[12846];
assign MEM[25444] = MEM[12623] + MEM[13639];
assign MEM[25445] = MEM[12627] + MEM[12987];
assign MEM[25446] = MEM[12632] + MEM[15368];
assign MEM[25447] = MEM[12635] + MEM[14495];
assign MEM[25448] = MEM[12636] + MEM[16915];
assign MEM[25449] = MEM[12637] + MEM[13128];
assign MEM[25450] = MEM[12639] + MEM[16460];
assign MEM[25451] = MEM[12640] + MEM[13124];
assign MEM[25452] = MEM[12647] + MEM[13501];
assign MEM[25453] = MEM[12648] + MEM[13365];
assign MEM[25454] = MEM[12651] + MEM[13645];
assign MEM[25455] = MEM[12653] + MEM[14427];
assign MEM[25456] = MEM[12654] + MEM[12895];
assign MEM[25457] = MEM[12655] + MEM[13050];
assign MEM[25458] = MEM[12658] + MEM[13683];
assign MEM[25459] = MEM[12665] + MEM[13923];
assign MEM[25460] = MEM[12669] + MEM[14311];
assign MEM[25461] = MEM[12673] + MEM[13563];
assign MEM[25462] = MEM[12675] + MEM[15011];
assign MEM[25463] = MEM[12677] + MEM[13481];
assign MEM[25464] = MEM[12679] + MEM[13243];
assign MEM[25465] = MEM[12680] + MEM[12769];
assign MEM[25466] = MEM[12681] + MEM[14875];
assign MEM[25467] = MEM[12683] + MEM[13127];
assign MEM[25468] = MEM[12684] + MEM[12808];
assign MEM[25469] = MEM[12687] + MEM[15802];
assign MEM[25470] = MEM[12690] + MEM[15180];
assign MEM[25471] = MEM[12691] + MEM[13724];
assign MEM[25472] = MEM[12696] + MEM[12858];
assign MEM[25473] = MEM[12698] + MEM[15164];
assign MEM[25474] = MEM[12702] + MEM[13181];
assign MEM[25475] = MEM[12703] + MEM[15504];
assign MEM[25476] = MEM[12706] + MEM[13880];
assign MEM[25477] = MEM[12712] + MEM[15392];
assign MEM[25478] = MEM[12713] + MEM[13774];
assign MEM[25479] = MEM[12716] + MEM[13402];
assign MEM[25480] = MEM[12717] + MEM[13859];
assign MEM[25481] = MEM[12719] + MEM[12870];
assign MEM[25482] = MEM[12721] + MEM[14612];
assign MEM[25483] = MEM[12723] + MEM[12973];
assign MEM[25484] = MEM[12724] + MEM[16605];
assign MEM[25485] = MEM[12725] + MEM[13743];
assign MEM[25486] = MEM[12726] + MEM[14292];
assign MEM[25487] = MEM[12728] + MEM[13191];
assign MEM[25488] = MEM[12731] + MEM[13857];
assign MEM[25489] = MEM[12740] + MEM[14064];
assign MEM[25490] = MEM[12742] + MEM[16018];
assign MEM[25491] = MEM[12744] + MEM[13870];
assign MEM[25492] = MEM[12745] + MEM[16284];
assign MEM[25493] = MEM[12747] + MEM[13908];
assign MEM[25494] = MEM[12753] + MEM[12925];
assign MEM[25495] = MEM[12754] + MEM[13200];
assign MEM[25496] = MEM[12756] + MEM[12783];
assign MEM[25497] = MEM[12759] + MEM[15381];
assign MEM[25498] = MEM[12764] + MEM[13247];
assign MEM[25499] = MEM[12770] + MEM[13482];
assign MEM[25500] = MEM[12771] + MEM[13409];
assign MEM[25501] = MEM[12778] + MEM[15006];
assign MEM[25502] = MEM[12779] + MEM[17518];
assign MEM[25503] = MEM[12781] + MEM[13710];
assign MEM[25504] = MEM[12782] + MEM[14999];
assign MEM[25505] = MEM[12787] + MEM[17218];
assign MEM[25506] = MEM[12788] + MEM[12871];
assign MEM[25507] = MEM[12789] + MEM[14952];
assign MEM[25508] = MEM[12792] + MEM[13814];
assign MEM[25509] = MEM[12797] + MEM[13960];
assign MEM[25510] = MEM[12798] + MEM[18096];
assign MEM[25511] = MEM[12800] + MEM[13626];
assign MEM[25512] = MEM[12801] + MEM[13519];
assign MEM[25513] = MEM[12802] + MEM[13871];
assign MEM[25514] = MEM[12803] + MEM[15787];
assign MEM[25515] = MEM[12806] + MEM[14372];
assign MEM[25516] = MEM[12809] + MEM[13242];
assign MEM[25517] = MEM[12814] + MEM[17136];
assign MEM[25518] = MEM[12822] + MEM[14992];
assign MEM[25519] = MEM[12824] + MEM[15804];
assign MEM[25520] = MEM[12825] + MEM[13499];
assign MEM[25521] = MEM[12826] + MEM[13095];
assign MEM[25522] = MEM[12829] + MEM[13727];
assign MEM[25523] = MEM[12830] + MEM[16097];
assign MEM[25524] = MEM[12834] + MEM[15047];
assign MEM[25525] = MEM[12836] + MEM[17778];
assign MEM[25526] = MEM[12837] + MEM[13332];
assign MEM[25527] = MEM[12839] + MEM[16268];
assign MEM[25528] = MEM[12841] + MEM[14206];
assign MEM[25529] = MEM[12843] + MEM[13604];
assign MEM[25530] = MEM[12845] + MEM[16847];
assign MEM[25531] = MEM[12848] + MEM[14435];
assign MEM[25532] = MEM[12851] + MEM[14406];
assign MEM[25533] = MEM[12859] + MEM[13763];
assign MEM[25534] = MEM[12864] + MEM[16796];
assign MEM[25535] = MEM[12865] + MEM[12992];
assign MEM[25536] = MEM[12866] + MEM[13715];
assign MEM[25537] = MEM[12867] + MEM[14561];
assign MEM[25538] = MEM[12872] + MEM[13199];
assign MEM[25539] = MEM[12875] + MEM[14788];
assign MEM[25540] = MEM[12876] + MEM[13811];
assign MEM[25541] = MEM[12880] + MEM[16602];
assign MEM[25542] = MEM[12881] + MEM[15050];
assign MEM[25543] = MEM[12883] + MEM[13596];
assign MEM[25544] = MEM[12890] + MEM[13812];
assign MEM[25545] = MEM[12891] + MEM[15962];
assign MEM[25546] = MEM[12892] + MEM[13764];
assign MEM[25547] = MEM[12894] + MEM[14218];
assign MEM[25548] = MEM[12896] + MEM[13698];
assign MEM[25549] = MEM[12901] + MEM[12957];
assign MEM[25550] = MEM[12906] + MEM[13368];
assign MEM[25551] = MEM[12910] + MEM[14076];
assign MEM[25552] = MEM[12911] + MEM[13676];
assign MEM[25553] = MEM[12912] + MEM[14942];
assign MEM[25554] = MEM[12913] + MEM[13391];
assign MEM[25555] = MEM[12914] + MEM[14358];
assign MEM[25556] = MEM[12918] + MEM[13362];
assign MEM[25557] = MEM[12919] + MEM[15994];
assign MEM[25558] = MEM[12920] + MEM[13731];
assign MEM[25559] = MEM[12922] + MEM[13215];
assign MEM[25560] = MEM[12923] + MEM[13188];
assign MEM[25561] = MEM[12924] + MEM[16561];
assign MEM[25562] = MEM[12926] + MEM[15343];
assign MEM[25563] = MEM[12928] + MEM[13237];
assign MEM[25564] = MEM[12933] + MEM[13121];
assign MEM[25565] = MEM[12934] + MEM[13788];
assign MEM[25566] = MEM[12940] + MEM[15116];
assign MEM[25567] = MEM[12943] + MEM[13492];
assign MEM[25568] = MEM[12944] + MEM[15254];
assign MEM[25569] = MEM[12946] + MEM[14881];
assign MEM[25570] = MEM[12947] + MEM[15242];
assign MEM[25571] = MEM[12951] + MEM[16258];
assign MEM[25572] = MEM[12952] + MEM[13538];
assign MEM[25573] = MEM[12954] + MEM[13571];
assign MEM[25574] = MEM[12955] + MEM[12994];
assign MEM[25575] = MEM[12958] + MEM[14148];
assign MEM[25576] = MEM[12959] + MEM[13278];
assign MEM[25577] = MEM[12960] + MEM[15868];
assign MEM[25578] = MEM[12964] + MEM[17526];
assign MEM[25579] = MEM[12967] + MEM[13406];
assign MEM[25580] = MEM[12974] + MEM[14642];
assign MEM[25581] = MEM[12975] + MEM[15617];
assign MEM[25582] = MEM[12980] + MEM[14674];
assign MEM[25583] = MEM[12981] + MEM[13893];
assign MEM[25584] = MEM[12990] + MEM[15429];
assign MEM[25585] = MEM[12995] + MEM[13742];
assign MEM[25586] = MEM[12996] + MEM[16493];
assign MEM[25587] = MEM[12998] + MEM[16552];
assign MEM[25588] = MEM[13001] + MEM[14317];
assign MEM[25589] = MEM[13003] + MEM[13468];
assign MEM[25590] = MEM[13008] + MEM[13105];
assign MEM[25591] = MEM[13010] + MEM[13671];
assign MEM[25592] = MEM[13011] + MEM[15841];
assign MEM[25593] = MEM[13013] + MEM[13163];
assign MEM[25594] = MEM[13016] + MEM[13030];
assign MEM[25595] = MEM[13018] + MEM[13785];
assign MEM[25596] = MEM[13026] + MEM[13465];
assign MEM[25597] = MEM[13027] + MEM[13077];
assign MEM[25598] = MEM[13031] + MEM[14294];
assign MEM[25599] = MEM[13033] + MEM[13062];
assign MEM[25600] = MEM[13034] + MEM[14474];
assign MEM[25601] = MEM[13035] + MEM[13227];
assign MEM[25602] = MEM[13037] + MEM[13713];
assign MEM[25603] = MEM[13038] + MEM[15531];
assign MEM[25604] = MEM[13039] + MEM[13319];
assign MEM[25605] = MEM[13043] + MEM[13600];
assign MEM[25606] = MEM[13049] + MEM[14763];
assign MEM[25607] = MEM[13051] + MEM[15512];
assign MEM[25608] = MEM[13052] + MEM[15364];
assign MEM[25609] = MEM[13056] + MEM[13544];
assign MEM[25610] = MEM[13061] + MEM[13898];
assign MEM[25611] = MEM[13063] + MEM[14058];
assign MEM[25612] = MEM[13065] + MEM[13285];
assign MEM[25613] = MEM[13069] + MEM[13490];
assign MEM[25614] = MEM[13071] + MEM[15502];
assign MEM[25615] = MEM[13073] + MEM[13196];
assign MEM[25616] = MEM[13075] + MEM[14476];
assign MEM[25617] = MEM[13078] + MEM[16779];
assign MEM[25618] = MEM[13081] + MEM[13096];
assign MEM[25619] = MEM[13082] + MEM[13432];
assign MEM[25620] = MEM[13084] + MEM[13991];
assign MEM[25621] = MEM[13089] + MEM[13286];
assign MEM[25622] = MEM[13091] + MEM[17024];
assign MEM[25623] = MEM[13097] + MEM[13145];
assign MEM[25624] = MEM[13098] + MEM[13565];
assign MEM[25625] = MEM[13100] + MEM[15340];
assign MEM[25626] = MEM[13101] + MEM[14108];
assign MEM[25627] = MEM[13103] + MEM[16504];
assign MEM[25628] = MEM[13106] + MEM[15371];
assign MEM[25629] = MEM[13109] + MEM[13295];
assign MEM[25630] = MEM[13114] + MEM[13894];
assign MEM[25631] = MEM[13118] + MEM[15999];
assign MEM[25632] = MEM[13120] + MEM[17017];
assign MEM[25633] = MEM[13123] + MEM[14267];
assign MEM[25634] = MEM[13126] + MEM[14086];
assign MEM[25635] = MEM[13130] + MEM[15562];
assign MEM[25636] = MEM[13132] + MEM[14819];
assign MEM[25637] = MEM[13136] + MEM[14047];
assign MEM[25638] = MEM[13138] + MEM[13558];
assign MEM[25639] = MEM[13139] + MEM[14194];
assign MEM[25640] = MEM[13141] + MEM[13906];
assign MEM[25641] = MEM[13142] + MEM[17122];
assign MEM[25642] = MEM[13143] + MEM[13386];
assign MEM[25643] = MEM[13148] + MEM[13545];
assign MEM[25644] = MEM[13152] + MEM[13364];
assign MEM[25645] = MEM[13157] + MEM[13315];
assign MEM[25646] = MEM[13158] + MEM[13791];
assign MEM[25647] = MEM[13162] + MEM[13622];
assign MEM[25648] = MEM[13173] + MEM[13178];
assign MEM[25649] = MEM[13175] + MEM[14025];
assign MEM[25650] = MEM[13177] + MEM[13616];
assign MEM[25651] = MEM[13180] + MEM[13310];
assign MEM[25652] = MEM[13187] + MEM[17290];
assign MEM[25653] = MEM[13190] + MEM[13588];
assign MEM[25654] = MEM[13192] + MEM[15932];
assign MEM[25655] = MEM[13193] + MEM[13516];
assign MEM[25656] = MEM[13205] + MEM[15692];
assign MEM[25657] = MEM[13207] + MEM[14011];
assign MEM[25658] = MEM[13210] + MEM[13621];
assign MEM[25659] = MEM[13211] + MEM[15167];
assign MEM[25660] = MEM[13217] + MEM[13714];
assign MEM[25661] = MEM[13219] + MEM[15354];
assign MEM[25662] = MEM[13220] + MEM[13668];
assign MEM[25663] = MEM[13224] + MEM[16196];
assign MEM[25664] = MEM[13226] + MEM[13307];
assign MEM[25665] = MEM[13231] + MEM[14134];
assign MEM[25666] = MEM[13232] + MEM[13598];
assign MEM[25667] = MEM[13235] + MEM[14455];
assign MEM[25668] = MEM[13245] + MEM[13434];
assign MEM[25669] = MEM[13248] + MEM[13826];
assign MEM[25670] = MEM[13249] + MEM[13273];
assign MEM[25671] = MEM[13251] + MEM[13360];
assign MEM[25672] = MEM[13252] + MEM[13524];
assign MEM[25673] = MEM[13256] + MEM[13341];
assign MEM[25674] = MEM[13258] + MEM[14809];
assign MEM[25675] = MEM[13259] + MEM[13268];
assign MEM[25676] = MEM[13264] + MEM[13407];
assign MEM[25677] = MEM[13269] + MEM[18047];
assign MEM[25678] = MEM[13276] + MEM[14338];
assign MEM[25679] = MEM[13284] + MEM[14356];
assign MEM[25680] = MEM[13288] + MEM[15326];
assign MEM[25681] = MEM[13290] + MEM[13863];
assign MEM[25682] = MEM[13292] + MEM[13578];
assign MEM[25683] = MEM[13294] + MEM[13564];
assign MEM[25684] = MEM[13296] + MEM[13822];
assign MEM[25685] = MEM[13297] + MEM[14753];
assign MEM[25686] = MEM[13298] + MEM[17298];
assign MEM[25687] = MEM[13299] + MEM[13934];
assign MEM[25688] = MEM[13304] + MEM[14123];
assign MEM[25689] = MEM[13305] + MEM[13720];
assign MEM[25690] = MEM[13308] + MEM[16624];
assign MEM[25691] = MEM[13311] + MEM[13560];
assign MEM[25692] = MEM[13313] + MEM[13507];
assign MEM[25693] = MEM[13314] + MEM[13705];
assign MEM[25694] = MEM[13318] + MEM[16008];
assign MEM[25695] = MEM[13324] + MEM[13670];
assign MEM[25696] = MEM[13325] + MEM[13531];
assign MEM[25697] = MEM[13326] + MEM[14070];
assign MEM[25698] = MEM[13327] + MEM[13421];
assign MEM[25699] = MEM[13328] + MEM[13660];
assign MEM[25700] = MEM[13329] + MEM[13597];
assign MEM[25701] = MEM[13331] + MEM[13846];
assign MEM[25702] = MEM[13333] + MEM[15143];
assign MEM[25703] = MEM[13334] + MEM[14769];
assign MEM[25704] = MEM[13337] + MEM[13393];
assign MEM[25705] = MEM[13339] + MEM[14071];
assign MEM[25706] = MEM[13340] + MEM[17201];
assign MEM[25707] = MEM[13344] + MEM[15571];
assign MEM[25708] = MEM[13346] + MEM[14986];
assign MEM[25709] = MEM[13347] + MEM[17383];
assign MEM[25710] = MEM[13354] + MEM[13982];
assign MEM[25711] = MEM[13355] + MEM[14561];
assign MEM[25712] = MEM[13361] + MEM[15064];
assign MEM[25713] = MEM[13366] + MEM[13630];
assign MEM[25714] = MEM[13369] + MEM[15785];
assign MEM[25715] = MEM[13371] + MEM[13380];
assign MEM[25716] = MEM[13374] + MEM[13976];
assign MEM[25717] = MEM[13378] + MEM[13431];
assign MEM[25718] = MEM[13382] + MEM[20740];
assign MEM[25719] = MEM[13389] + MEM[13940];
assign MEM[25720] = MEM[13396] + MEM[14743];
assign MEM[25721] = MEM[13399] + MEM[14381];
assign MEM[25722] = MEM[13403] + MEM[14887];
assign MEM[25723] = MEM[13408] + MEM[14823];
assign MEM[25724] = MEM[13411] + MEM[15179];
assign MEM[25725] = MEM[13413] + MEM[15144];
assign MEM[25726] = MEM[13416] + MEM[14695];
assign MEM[25727] = MEM[13427] + MEM[15053];
assign MEM[25728] = MEM[13430] + MEM[18793];
assign MEM[25729] = MEM[13433] + MEM[15871];
assign MEM[25730] = MEM[13436] + MEM[13551];
assign MEM[25731] = MEM[13437] + MEM[14691];
assign MEM[25732] = MEM[13438] + MEM[13704];
assign MEM[25733] = MEM[13439] + MEM[13480];
assign MEM[25734] = MEM[13443] + MEM[15572];
assign MEM[25735] = MEM[13444] + MEM[13917];
assign MEM[25736] = MEM[13448] + MEM[15691];
assign MEM[25737] = MEM[13451] + MEM[13978];
assign MEM[25738] = MEM[13454] + MEM[20179];
assign MEM[25739] = MEM[13458] + MEM[14762];
assign MEM[25740] = MEM[13459] + MEM[15867];
assign MEM[25741] = MEM[13460] + MEM[15938];
assign MEM[25742] = MEM[13462] + MEM[13913];
assign MEM[25743] = MEM[13464] + MEM[15117];
assign MEM[25744] = MEM[13467] + MEM[15317];
assign MEM[25745] = MEM[13470] + MEM[15461];
assign MEM[25746] = MEM[13472] + MEM[13691];
assign MEM[25747] = MEM[13475] + MEM[13827];
assign MEM[25748] = MEM[13477] + MEM[13837];
assign MEM[25749] = MEM[13484] + MEM[15372];
assign MEM[25750] = MEM[13485] + MEM[14569];
assign MEM[25751] = MEM[13486] + MEM[14575];
assign MEM[25752] = MEM[13491] + MEM[14003];
assign MEM[25753] = MEM[13494] + MEM[14775];
assign MEM[25754] = MEM[13502] + MEM[14844];
assign MEM[25755] = MEM[13504] + MEM[14149];
assign MEM[25756] = MEM[13505] + MEM[15273];
assign MEM[25757] = MEM[13511] + MEM[13534];
assign MEM[25758] = MEM[13517] + MEM[16630];
assign MEM[25759] = MEM[13518] + MEM[15513];
assign MEM[25760] = MEM[13521] + MEM[16634];
assign MEM[25761] = MEM[13525] + MEM[13627];
assign MEM[25762] = MEM[13526] + MEM[15438];
assign MEM[25763] = MEM[13528] + MEM[13675];
assign MEM[25764] = MEM[13529] + MEM[13610];
assign MEM[25765] = MEM[13530] + MEM[13754];
assign MEM[25766] = MEM[13535] + MEM[15237];
assign MEM[25767] = MEM[13537] + MEM[17653];
assign MEM[25768] = MEM[13540] + MEM[18228];
assign MEM[25769] = MEM[13548] + MEM[13782];
assign MEM[25770] = MEM[13549] + MEM[18281];
assign MEM[25771] = MEM[13550] + MEM[13568];
assign MEM[25772] = MEM[13554] + MEM[16200];
assign MEM[25773] = MEM[13555] + MEM[13695];
assign MEM[25774] = MEM[13556] + MEM[13875];
assign MEM[25775] = MEM[13562] + MEM[15091];
assign MEM[25776] = MEM[13566] + MEM[16170];
assign MEM[25777] = MEM[13567] + MEM[13615];
assign MEM[25778] = MEM[13570] + MEM[13820];
assign MEM[25779] = MEM[13575] + MEM[14984];
assign MEM[25780] = MEM[13576] + MEM[14125];
assign MEM[25781] = MEM[13577] + MEM[16171];
assign MEM[25782] = MEM[13579] + MEM[14164];
assign MEM[25783] = MEM[13582] + MEM[14043];
assign MEM[25784] = MEM[13584] + MEM[14050];
assign MEM[25785] = MEM[13585] + MEM[15761];
assign MEM[25786] = MEM[13590] + MEM[13650];
assign MEM[25787] = MEM[13591] + MEM[16478];
assign MEM[25788] = MEM[13592] + MEM[13749];
assign MEM[25789] = MEM[13593] + MEM[15090];
assign MEM[25790] = MEM[13599] + MEM[14307];
assign MEM[25791] = MEM[13601] + MEM[13919];
assign MEM[25792] = MEM[13606] + MEM[14426];
assign MEM[25793] = MEM[13607] + MEM[18495];
assign MEM[25794] = MEM[13611] + MEM[15844];
assign MEM[25795] = MEM[13613] + MEM[15311];
assign MEM[25796] = MEM[13614] + MEM[13885];
assign MEM[25797] = MEM[13618] + MEM[14262];
assign MEM[25798] = MEM[13619] + MEM[14331];
assign MEM[25799] = MEM[13625] + MEM[13771];
assign MEM[25800] = MEM[13628] + MEM[14567];
assign MEM[25801] = MEM[13629] + MEM[14859];
assign MEM[25802] = MEM[13631] + MEM[16163];
assign MEM[25803] = MEM[13643] + MEM[13707];
assign MEM[25804] = MEM[13646] + MEM[15735];
assign MEM[25805] = MEM[13647] + MEM[14822];
assign MEM[25806] = MEM[13654] + MEM[14077];
assign MEM[25807] = MEM[13656] + MEM[14126];
assign MEM[25808] = MEM[13661] + MEM[13673];
assign MEM[25809] = MEM[13663] + MEM[13730];
assign MEM[25810] = MEM[13664] + MEM[15963];
assign MEM[25811] = MEM[13669] + MEM[14675];
assign MEM[25812] = MEM[13682] + MEM[13794];
assign MEM[25813] = MEM[13684] + MEM[13942];
assign MEM[25814] = MEM[13689] + MEM[14083];
assign MEM[25815] = MEM[13692] + MEM[14729];
assign MEM[25816] = MEM[13693] + MEM[14721];
assign MEM[25817] = MEM[13696] + MEM[15257];
assign MEM[25818] = MEM[13708] + MEM[15317];
assign MEM[25819] = MEM[13709] + MEM[13747];
assign MEM[25820] = MEM[13712] + MEM[14296];
assign MEM[25821] = MEM[13716] + MEM[18784];
assign MEM[25822] = MEM[13717] + MEM[15332];
assign MEM[25823] = MEM[13718] + MEM[14145];
assign MEM[25824] = MEM[13722] + MEM[13735];
assign MEM[25825] = MEM[13723] + MEM[15882];
assign MEM[25826] = MEM[13726] + MEM[14907];
assign MEM[25827] = MEM[13728] + MEM[17013];
assign MEM[25828] = MEM[13732] + MEM[17054];
assign MEM[25829] = MEM[13733] + MEM[13900];
assign MEM[25830] = MEM[13734] + MEM[15516];
assign MEM[25831] = MEM[13736] + MEM[15673];
assign MEM[25832] = MEM[13737] + MEM[14416];
assign MEM[25833] = MEM[13738] + MEM[15430];
assign MEM[25834] = MEM[13740] + MEM[14056];
assign MEM[25835] = MEM[13741] + MEM[15820];
assign MEM[25836] = MEM[13744] + MEM[16061];
assign MEM[25837] = MEM[13750] + MEM[15044];
assign MEM[25838] = MEM[13752] + MEM[14171];
assign MEM[25839] = MEM[13761] + MEM[13925];
assign MEM[25840] = MEM[13762] + MEM[14005];
assign MEM[25841] = MEM[13765] + MEM[14429];
assign MEM[25842] = MEM[13766] + MEM[14439];
assign MEM[25843] = MEM[13767] + MEM[14429];
assign MEM[25844] = MEM[13768] + MEM[16233];
assign MEM[25845] = MEM[13773] + MEM[13789];
assign MEM[25846] = MEM[13778] + MEM[14039];
assign MEM[25847] = MEM[13783] + MEM[14390];
assign MEM[25848] = MEM[13784] + MEM[16253];
assign MEM[25849] = MEM[13786] + MEM[18473];
assign MEM[25850] = MEM[13792] + MEM[15804];
assign MEM[25851] = MEM[13796] + MEM[15948];
assign MEM[25852] = MEM[13798] + MEM[16040];
assign MEM[25853] = MEM[13801] + MEM[18073];
assign MEM[25854] = MEM[13802] + MEM[15882];
assign MEM[25855] = MEM[13804] + MEM[16603];
assign MEM[25856] = MEM[13810] + MEM[14781];
assign MEM[25857] = MEM[13813] + MEM[15422];
assign MEM[25858] = MEM[13815] + MEM[16207];
assign MEM[25859] = MEM[13817] + MEM[14669];
assign MEM[25860] = MEM[13818] + MEM[15503];
assign MEM[25861] = MEM[13819] + MEM[14136];
assign MEM[25862] = MEM[13827] + MEM[16189];
assign MEM[25863] = MEM[13828] + MEM[15609];
assign MEM[25864] = MEM[13830] + MEM[14796];
assign MEM[25865] = MEM[13831] + MEM[14040];
assign MEM[25866] = MEM[13832] + MEM[14127];
assign MEM[25867] = MEM[13833] + MEM[15601];
assign MEM[25868] = MEM[13834] + MEM[15000];
assign MEM[25869] = MEM[13836] + MEM[15770];
assign MEM[25870] = MEM[13838] + MEM[14639];
assign MEM[25871] = MEM[13840] + MEM[14015];
assign MEM[25872] = MEM[13841] + MEM[14334];
assign MEM[25873] = MEM[13842] + MEM[16926];
assign MEM[25874] = MEM[13843] + MEM[14242];
assign MEM[25875] = MEM[13845] + MEM[17273];
assign MEM[25876] = MEM[13847] + MEM[17750];
assign MEM[25877] = MEM[13850] + MEM[16525];
assign MEM[25878] = MEM[13851] + MEM[16541];
assign MEM[25879] = MEM[13852] + MEM[14412];
assign MEM[25880] = MEM[13853] + MEM[14072];
assign MEM[25881] = MEM[13854] + MEM[14586];
assign MEM[25882] = MEM[13855] + MEM[14723];
assign MEM[25883] = MEM[13856] + MEM[16094];
assign MEM[25884] = MEM[13858] + MEM[15587];
assign MEM[25885] = MEM[13860] + MEM[16137];
assign MEM[25886] = MEM[13861] + MEM[15853];
assign MEM[25887] = MEM[13862] + MEM[16912];
assign MEM[25888] = MEM[13864] + MEM[14605];
assign MEM[25889] = MEM[13867] + MEM[14221];
assign MEM[25890] = MEM[13868] + MEM[15995];
assign MEM[25891] = MEM[13869] + MEM[14314];
assign MEM[25892] = MEM[13872] + MEM[14589];
assign MEM[25893] = MEM[13873] + MEM[14526];
assign MEM[25894] = MEM[13876] + MEM[15375];
assign MEM[25895] = MEM[13877] + MEM[13910];
assign MEM[25896] = MEM[13878] + MEM[14804];
assign MEM[25897] = MEM[13879] + MEM[14304];
assign MEM[25898] = MEM[13881] + MEM[15816];
assign MEM[25899] = MEM[13882] + MEM[15776];
assign MEM[25900] = MEM[13883] + MEM[18185];
assign MEM[25901] = MEM[13884] + MEM[16163];
assign MEM[25902] = MEM[13886] + MEM[14176];
assign MEM[25903] = MEM[13888] + MEM[15924];
assign MEM[25904] = MEM[13889] + MEM[13928];
assign MEM[25905] = MEM[13891] + MEM[15289];
assign MEM[25906] = MEM[13892] + MEM[15875];
assign MEM[25907] = MEM[13895] + MEM[14073];
assign MEM[25908] = MEM[13896] + MEM[17675];
assign MEM[25909] = MEM[13901] + MEM[15008];
assign MEM[25910] = MEM[13902] + MEM[15126];
assign MEM[25911] = MEM[13903] + MEM[15284];
assign MEM[25912] = MEM[13904] + MEM[16656];
assign MEM[25913] = MEM[13905] + MEM[15356];
assign MEM[25914] = MEM[13907] + MEM[16403];
assign MEM[25915] = MEM[13911] + MEM[15228];
assign MEM[25916] = MEM[13912] + MEM[14932];
assign MEM[25917] = MEM[13914] + MEM[15724];
assign MEM[25918] = MEM[13915] + MEM[16059];
assign MEM[25919] = MEM[13918] + MEM[17019];
assign MEM[25920] = MEM[13922] + MEM[15771];
assign MEM[25921] = MEM[13924] + MEM[14022];
assign MEM[25922] = MEM[13926] + MEM[17032];
assign MEM[25923] = MEM[13927] + MEM[14890];
assign MEM[25924] = MEM[13930] + MEM[14891];
assign MEM[25925] = MEM[13931] + MEM[14798];
assign MEM[25926] = MEM[13933] + MEM[16636];
assign MEM[25927] = MEM[13935] + MEM[14131];
assign MEM[25928] = MEM[13936] + MEM[14316];
assign MEM[25929] = MEM[13937] + MEM[14567];
assign MEM[25930] = MEM[13941] + MEM[16195];
assign MEM[25931] = MEM[13943] + MEM[17429];
assign MEM[25932] = MEM[13944] + MEM[17554];
assign MEM[25933] = MEM[13945] + MEM[15186];
assign MEM[25934] = MEM[13946] + MEM[14065];
assign MEM[25935] = MEM[13947] + MEM[15576];
assign MEM[25936] = MEM[13948] + MEM[16273];
assign MEM[25937] = MEM[13949] + MEM[14583];
assign MEM[25938] = MEM[13950] + MEM[16401];
assign MEM[25939] = MEM[13951] + MEM[14000];
assign MEM[25940] = MEM[13952] + MEM[14254];
assign MEM[25941] = MEM[13953] + MEM[14523];
assign MEM[25942] = MEM[13955] + MEM[15449];
assign MEM[25943] = MEM[13956] + MEM[17897];
assign MEM[25944] = MEM[13957] + MEM[14220];
assign MEM[25945] = MEM[13958] + MEM[16025];
assign MEM[25946] = MEM[13959] + MEM[16868];
assign MEM[25947] = MEM[13961] + MEM[15640];
assign MEM[25948] = MEM[13962] + MEM[14890];
assign MEM[25949] = MEM[13964] + MEM[16287];
assign MEM[25950] = MEM[13966] + MEM[14030];
assign MEM[25951] = MEM[13967] + MEM[15389];
assign MEM[25952] = MEM[13969] + MEM[18505];
assign MEM[25953] = MEM[13970] + MEM[14172];
assign MEM[25954] = MEM[13971] + MEM[15635];
assign MEM[25955] = MEM[13972] + MEM[16046];
assign MEM[25956] = MEM[13974] + MEM[14054];
assign MEM[25957] = MEM[13975] + MEM[14735];
assign MEM[25958] = MEM[13977] + MEM[16211];
assign MEM[25959] = MEM[13979] + MEM[17007];
assign MEM[25960] = MEM[13980] + MEM[17705];
assign MEM[25961] = MEM[13981] + MEM[16165];
assign MEM[25962] = MEM[13984] + MEM[19017];
assign MEM[25963] = MEM[13985] + MEM[15021];
assign MEM[25964] = MEM[13986] + MEM[15043];
assign MEM[25965] = MEM[13987] + MEM[15927];
assign MEM[25966] = MEM[13988] + MEM[15131];
assign MEM[25967] = MEM[13989] + MEM[16738];
assign MEM[25968] = MEM[13992] + MEM[15965];
assign MEM[25969] = MEM[13993] + MEM[16390];
assign MEM[25970] = MEM[13994] + MEM[14130];
assign MEM[25971] = MEM[13995] + MEM[15342];
assign MEM[25972] = MEM[13996] + MEM[15081];
assign MEM[25973] = MEM[13997] + MEM[14256];
assign MEM[25974] = MEM[13999] + MEM[14904];
assign MEM[25975] = MEM[14001] + MEM[14524];
assign MEM[25976] = MEM[14002] + MEM[17632];
assign MEM[25977] = MEM[14004] + MEM[16282];
assign MEM[25978] = MEM[14006] + MEM[15808];
assign MEM[25979] = MEM[14007] + MEM[14719];
assign MEM[25980] = MEM[14010] + MEM[14636];
assign MEM[25981] = MEM[14012] + MEM[14705];
assign MEM[25982] = MEM[14014] + MEM[14154];
assign MEM[25983] = MEM[14016] + MEM[15515];
assign MEM[25984] = MEM[14018] + MEM[16987];
assign MEM[25985] = MEM[14020] + MEM[14413];
assign MEM[25986] = MEM[14021] + MEM[14906];
assign MEM[25987] = MEM[14027] + MEM[15634];
assign MEM[25988] = MEM[14028] + MEM[14693];
assign MEM[25989] = MEM[14029] + MEM[15666];
assign MEM[25990] = MEM[14031] + MEM[14588];
assign MEM[25991] = MEM[14032] + MEM[15146];
assign MEM[25992] = MEM[14033] + MEM[14922];
assign MEM[25993] = MEM[14034] + MEM[14150];
assign MEM[25994] = MEM[14035] + MEM[15074];
assign MEM[25995] = MEM[14036] + MEM[18625];
assign MEM[25996] = MEM[14037] + MEM[16958];
assign MEM[25997] = MEM[14038] + MEM[16317];
assign MEM[25998] = MEM[14045] + MEM[15670];
assign MEM[25999] = MEM[14051] + MEM[14556];
assign MEM[26000] = MEM[14052] + MEM[14959];
assign MEM[26001] = MEM[14053] + MEM[17093];
assign MEM[26002] = MEM[14055] + MEM[14530];
assign MEM[26003] = MEM[14057] + MEM[16686];
assign MEM[26004] = MEM[14059] + MEM[16691];
assign MEM[26005] = MEM[14060] + MEM[14882];
assign MEM[26006] = MEM[14061] + MEM[14184];
assign MEM[26007] = MEM[14062] + MEM[18336];
assign MEM[26008] = MEM[14063] + MEM[19416];
assign MEM[26009] = MEM[14066] + MEM[14988];
assign MEM[26010] = MEM[14067] + MEM[16777];
assign MEM[26011] = MEM[14068] + MEM[16740];
assign MEM[26012] = MEM[14074] + MEM[14434];
assign MEM[26013] = MEM[14081] + MEM[19125];
assign MEM[26014] = MEM[14085] + MEM[16126];
assign MEM[26015] = MEM[14087] + MEM[17422];
assign MEM[26016] = MEM[14088] + MEM[14279];
assign MEM[26017] = MEM[14089] + MEM[14544];
assign MEM[26018] = MEM[14090] + MEM[14623];
assign MEM[26019] = MEM[14091] + MEM[16518];
assign MEM[26020] = MEM[14092] + MEM[16192];
assign MEM[26021] = MEM[14093] + MEM[16028];
assign MEM[26022] = MEM[14094] + MEM[17427];
assign MEM[26023] = MEM[14098] + MEM[17853];
assign MEM[26024] = MEM[14099] + MEM[14814];
assign MEM[26025] = MEM[14101] + MEM[15321];
assign MEM[26026] = MEM[14102] + MEM[15286];
assign MEM[26027] = MEM[14103] + MEM[15968];
assign MEM[26028] = MEM[14105] + MEM[14575];
assign MEM[26029] = MEM[14107] + MEM[16301];
assign MEM[26030] = MEM[14109] + MEM[14509];
assign MEM[26031] = MEM[14110] + MEM[16185];
assign MEM[26032] = MEM[14111] + MEM[15080];
assign MEM[26033] = MEM[14113] + MEM[14361];
assign MEM[26034] = MEM[14114] + MEM[16221];
assign MEM[26035] = MEM[14115] + MEM[18104];
assign MEM[26036] = MEM[14116] + MEM[16612];
assign MEM[26037] = MEM[14118] + MEM[14580];
assign MEM[26038] = MEM[14119] + MEM[14724];
assign MEM[26039] = MEM[14121] + MEM[17056];
assign MEM[26040] = MEM[14122] + MEM[17125];
assign MEM[26041] = MEM[14124] + MEM[18716];
assign MEM[26042] = MEM[14128] + MEM[15897];
assign MEM[26043] = MEM[14129] + MEM[17428];
assign MEM[26044] = MEM[14132] + MEM[16764];
assign MEM[26045] = MEM[14133] + MEM[14470];
assign MEM[26046] = MEM[14135] + MEM[16170];
assign MEM[26047] = MEM[14137] + MEM[15269];
assign MEM[26048] = MEM[14138] + MEM[15645];
assign MEM[26049] = MEM[14139] + MEM[14513];
assign MEM[26050] = MEM[14140] + MEM[14541];
assign MEM[26051] = MEM[14142] + MEM[15402];
assign MEM[26052] = MEM[14143] + MEM[15607];
assign MEM[26053] = MEM[14146] + MEM[14595];
assign MEM[26054] = MEM[14151] + MEM[17029];
assign MEM[26055] = MEM[14153] + MEM[17326];
assign MEM[26056] = MEM[14155] + MEM[14811];
assign MEM[26057] = MEM[14156] + MEM[16031];
assign MEM[26058] = MEM[14157] + MEM[17473];
assign MEM[26059] = MEM[14159] + MEM[16287];
assign MEM[26060] = MEM[14160] + MEM[15240];
assign MEM[26061] = MEM[14161] + MEM[14969];
assign MEM[26062] = MEM[14162] + MEM[14204];
assign MEM[26063] = MEM[14163] + MEM[16013];
assign MEM[26064] = MEM[14165] + MEM[16228];
assign MEM[26065] = MEM[14166] + MEM[14271];
assign MEM[26066] = MEM[14168] + MEM[17917];
assign MEM[26067] = MEM[14169] + MEM[17483];
assign MEM[26068] = MEM[14170] + MEM[16181];
assign MEM[26069] = MEM[14173] + MEM[18771];
assign MEM[26070] = MEM[14174] + MEM[16701];
assign MEM[26071] = MEM[14177] + MEM[15377];
assign MEM[26072] = MEM[14179] + MEM[15471];
assign MEM[26073] = MEM[14180] + MEM[15136];
assign MEM[26074] = MEM[14181] + MEM[16442];
assign MEM[26075] = MEM[14182] + MEM[14211];
assign MEM[26076] = MEM[14183] + MEM[14185];
assign MEM[26077] = MEM[14186] + MEM[18581];
assign MEM[26078] = MEM[14187] + MEM[14698];
assign MEM[26079] = MEM[14188] + MEM[17065];
assign MEM[26080] = MEM[14189] + MEM[18545];
assign MEM[26081] = MEM[14190] + MEM[16723];
assign MEM[26082] = MEM[14191] + MEM[14401];
assign MEM[26083] = MEM[14192] + MEM[15007];
assign MEM[26084] = MEM[14193] + MEM[16049];
assign MEM[26085] = MEM[14195] + MEM[16872];
assign MEM[26086] = MEM[14196] + MEM[15062];
assign MEM[26087] = MEM[14197] + MEM[14202];
assign MEM[26088] = MEM[14198] + MEM[16733];
assign MEM[26089] = MEM[14199] + MEM[14658];
assign MEM[26090] = MEM[14200] + MEM[16563];
assign MEM[26091] = MEM[14201] + MEM[14607];
assign MEM[26092] = MEM[14203] + MEM[16865];
assign MEM[26093] = MEM[14209] + MEM[17045];
assign MEM[26094] = MEM[14212] + MEM[16422];
assign MEM[26095] = MEM[14213] + MEM[14378];
assign MEM[26096] = MEM[14214] + MEM[14465];
assign MEM[26097] = MEM[14219] + MEM[14252];
assign MEM[26098] = MEM[14222] + MEM[14324];
assign MEM[26099] = MEM[14223] + MEM[17053];
assign MEM[26100] = MEM[14225] + MEM[14532];
assign MEM[26101] = MEM[14226] + MEM[14278];
assign MEM[26102] = MEM[14228] + MEM[15262];
assign MEM[26103] = MEM[14229] + MEM[17826];
assign MEM[26104] = MEM[14230] + MEM[17642];
assign MEM[26105] = MEM[14232] + MEM[14877];
assign MEM[26106] = MEM[14233] + MEM[17738];
assign MEM[26107] = MEM[14234] + MEM[17474];
assign MEM[26108] = MEM[14236] + MEM[17423];
assign MEM[26109] = MEM[14237] + MEM[14490];
assign MEM[26110] = MEM[14239] + MEM[14418];
assign MEM[26111] = MEM[14240] + MEM[17561];
assign MEM[26112] = MEM[14241] + MEM[17506];
assign MEM[26113] = MEM[14246] + MEM[14977];
assign MEM[26114] = MEM[14247] + MEM[15702];
assign MEM[26115] = MEM[14248] + MEM[14367];
assign MEM[26116] = MEM[14249] + MEM[18260];
assign MEM[26117] = MEM[14250] + MEM[15097];
assign MEM[26118] = MEM[14251] + MEM[14460];
assign MEM[26119] = MEM[14255] + MEM[17618];
assign MEM[26120] = MEM[14257] + MEM[17730];
assign MEM[26121] = MEM[14261] + MEM[17943];
assign MEM[26122] = MEM[14264] + MEM[14951];
assign MEM[26123] = MEM[14265] + MEM[17510];
assign MEM[26124] = MEM[14266] + MEM[15381];
assign MEM[26125] = MEM[14268] + MEM[16638];
assign MEM[26126] = MEM[14269] + MEM[14980];
assign MEM[26127] = MEM[14270] + MEM[14430];
assign MEM[26128] = MEM[14272] + MEM[17262];
assign MEM[26129] = MEM[14274] + MEM[14989];
assign MEM[26130] = MEM[14275] + MEM[16695];
assign MEM[26131] = MEM[14276] + MEM[18002];
assign MEM[26132] = MEM[14277] + MEM[16521];
assign MEM[26133] = MEM[14278] + MEM[14614];
assign MEM[26134] = MEM[14280] + MEM[15951];
assign MEM[26135] = MEM[14281] + MEM[15445];
assign MEM[26136] = MEM[14282] + MEM[16138];
assign MEM[26137] = MEM[14283] + MEM[15974];
assign MEM[26138] = MEM[14285] + MEM[15441];
assign MEM[26139] = MEM[14288] + MEM[15484];
assign MEM[26140] = MEM[14289] + MEM[14759];
assign MEM[26141] = MEM[14290] + MEM[16954];
assign MEM[26142] = MEM[14291] + MEM[15208];
assign MEM[26143] = MEM[14293] + MEM[14504];
assign MEM[26144] = MEM[14295] + MEM[14487];
assign MEM[26145] = MEM[14297] + MEM[17615];
assign MEM[26146] = MEM[14299] + MEM[15774];
assign MEM[26147] = MEM[14300] + MEM[16864];
assign MEM[26148] = MEM[14301] + MEM[16989];
assign MEM[26149] = MEM[14302] + MEM[14857];
assign MEM[26150] = MEM[14303] + MEM[16402];
assign MEM[26151] = MEM[14305] + MEM[14944];
assign MEM[26152] = MEM[14306] + MEM[15235];
assign MEM[26153] = MEM[14309] + MEM[17082];
assign MEM[26154] = MEM[14312] + MEM[16961];
assign MEM[26155] = MEM[14313] + MEM[14998];
assign MEM[26156] = MEM[14318] + MEM[14899];
assign MEM[26157] = MEM[14319] + MEM[14838];
assign MEM[26158] = MEM[14320] + MEM[17641];
assign MEM[26159] = MEM[14321] + MEM[15646];
assign MEM[26160] = MEM[14322] + MEM[15876];
assign MEM[26161] = MEM[14323] + MEM[15983];
assign MEM[26162] = MEM[14325] + MEM[14330];
assign MEM[26163] = MEM[14326] + MEM[14382];
assign MEM[26164] = MEM[14327] + MEM[14344];
assign MEM[26165] = MEM[14328] + MEM[16585];
assign MEM[26166] = MEM[14329] + MEM[15587];
assign MEM[26167] = MEM[14332] + MEM[14791];
assign MEM[26168] = MEM[14333] + MEM[16317];
assign MEM[26169] = MEM[14339] + MEM[18613];
assign MEM[26170] = MEM[14340] + MEM[16565];
assign MEM[26171] = MEM[14341] + MEM[16579];
assign MEM[26172] = MEM[14343] + MEM[16166];
assign MEM[26173] = MEM[14345] + MEM[16368];
assign MEM[26174] = MEM[14347] + MEM[16614];
assign MEM[26175] = MEM[14348] + MEM[15159];
assign MEM[26176] = MEM[14349] + MEM[16759];
assign MEM[26177] = MEM[14350] + MEM[14919];
assign MEM[26178] = MEM[14351] + MEM[18492];
assign MEM[26179] = MEM[14352] + MEM[14739];
assign MEM[26180] = MEM[14353] + MEM[16338];
assign MEM[26181] = MEM[14354] + MEM[15437];
assign MEM[26182] = MEM[14357] + MEM[18184];
assign MEM[26183] = MEM[14359] + MEM[17639];
assign MEM[26184] = MEM[14360] + MEM[15716];
assign MEM[26185] = MEM[14362] + MEM[14794];
assign MEM[26186] = MEM[14364] + MEM[14990];
assign MEM[26187] = MEM[14365] + MEM[16175];
assign MEM[26188] = MEM[14368] + MEM[17956];
assign MEM[26189] = MEM[14369] + MEM[15024];
assign MEM[26190] = MEM[14370] + MEM[14847];
assign MEM[26191] = MEM[14371] + MEM[14507];
assign MEM[26192] = MEM[14373] + MEM[15233];
assign MEM[26193] = MEM[14375] + MEM[18116];
assign MEM[26194] = MEM[14376] + MEM[14621];
assign MEM[26195] = MEM[14380] + MEM[19788];
assign MEM[26196] = MEM[14383] + MEM[15606];
assign MEM[26197] = MEM[14386] + MEM[15591];
assign MEM[26198] = MEM[14388] + MEM[14865];
assign MEM[26199] = MEM[14391] + MEM[17646];
assign MEM[26200] = MEM[14392] + MEM[14670];
assign MEM[26201] = MEM[14393] + MEM[14808];
assign MEM[26202] = MEM[14394] + MEM[16790];
assign MEM[26203] = MEM[14395] + MEM[17588];
assign MEM[26204] = MEM[14396] + MEM[16422];
assign MEM[26205] = MEM[14397] + MEM[17676];
assign MEM[26206] = MEM[14398] + MEM[15780];
assign MEM[26207] = MEM[14400] + MEM[17197];
assign MEM[26208] = MEM[14402] + MEM[17051];
assign MEM[26209] = MEM[14403] + MEM[15598];
assign MEM[26210] = MEM[14404] + MEM[14853];
assign MEM[26211] = MEM[14405] + MEM[16627];
assign MEM[26212] = MEM[14407] + MEM[16711];
assign MEM[26213] = MEM[14410] + MEM[15390];
assign MEM[26214] = MEM[14411] + MEM[17364];
assign MEM[26215] = MEM[14414] + MEM[14750];
assign MEM[26216] = MEM[14415] + MEM[17558];
assign MEM[26217] = MEM[14419] + MEM[17519];
assign MEM[26218] = MEM[14420] + MEM[14577];
assign MEM[26219] = MEM[14421] + MEM[14643];
assign MEM[26220] = MEM[14422] + MEM[14746];
assign MEM[26221] = MEM[14423] + MEM[14917];
assign MEM[26222] = MEM[14424] + MEM[14581];
assign MEM[26223] = MEM[14425] + MEM[15929];
assign MEM[26224] = MEM[14431] + MEM[14961];
assign MEM[26225] = MEM[14432] + MEM[17812];
assign MEM[26226] = MEM[14433] + MEM[15432];
assign MEM[26227] = MEM[14436] + MEM[17596];
assign MEM[26228] = MEM[14437] + MEM[18322];
assign MEM[26229] = MEM[14438] + MEM[19485];
assign MEM[26230] = MEM[14440] + MEM[15762];
assign MEM[26231] = MEM[14441] + MEM[15691];
assign MEM[26232] = MEM[14442] + MEM[15674];
assign MEM[26233] = MEM[14443] + MEM[18055];
assign MEM[26234] = MEM[14445] + MEM[14736];
assign MEM[26235] = MEM[14446] + MEM[15243];
assign MEM[26236] = MEM[14447] + MEM[14731];
assign MEM[26237] = MEM[14448] + MEM[15555];
assign MEM[26238] = MEM[14450] + MEM[17279];
assign MEM[26239] = MEM[14451] + MEM[15819];
assign MEM[26240] = MEM[14452] + MEM[15123];
assign MEM[26241] = MEM[14454] + MEM[14913];
assign MEM[26242] = MEM[14457] + MEM[14629];
assign MEM[26243] = MEM[14458] + MEM[17566];
assign MEM[26244] = MEM[14459] + MEM[17104];
assign MEM[26245] = MEM[14461] + MEM[17552];
assign MEM[26246] = MEM[14462] + MEM[17688];
assign MEM[26247] = MEM[14463] + MEM[14560];
assign MEM[26248] = MEM[14466] + MEM[16499];
assign MEM[26249] = MEM[14467] + MEM[14749];
assign MEM[26250] = MEM[14468] + MEM[18356];
assign MEM[26251] = MEM[14469] + MEM[14542];
assign MEM[26252] = MEM[14471] + MEM[16531];
assign MEM[26253] = MEM[14472] + MEM[15984];
assign MEM[26254] = MEM[14473] + MEM[18382];
assign MEM[26255] = MEM[14475] + MEM[15910];
assign MEM[26256] = MEM[14477] + MEM[14975];
assign MEM[26257] = MEM[14478] + MEM[18796];
assign MEM[26258] = MEM[14479] + MEM[17286];
assign MEM[26259] = MEM[14480] + MEM[14529];
assign MEM[26260] = MEM[14481] + MEM[14535];
assign MEM[26261] = MEM[14482] + MEM[16547];
assign MEM[26262] = MEM[14483] + MEM[15056];
assign MEM[26263] = MEM[14484] + MEM[15369];
assign MEM[26264] = MEM[14485] + MEM[15570];
assign MEM[26265] = MEM[14486] + MEM[15807];
assign MEM[26266] = MEM[14488] + MEM[14845];
assign MEM[26267] = MEM[14489] + MEM[16073];
assign MEM[26268] = MEM[14491] + MEM[14640];
assign MEM[26269] = MEM[14494] + MEM[14832];
assign MEM[26270] = MEM[14496] + MEM[17050];
assign MEM[26271] = MEM[14498] + MEM[15987];
assign MEM[26272] = MEM[14499] + MEM[15092];
assign MEM[26273] = MEM[14500] + MEM[14820];
assign MEM[26274] = MEM[14502] + MEM[17512];
assign MEM[26275] = MEM[14505] + MEM[14768];
assign MEM[26276] = MEM[14506] + MEM[15218];
assign MEM[26277] = MEM[14508] + MEM[15017];
assign MEM[26278] = MEM[14510] + MEM[16908];
assign MEM[26279] = MEM[14511] + MEM[17725];
assign MEM[26280] = MEM[14512] + MEM[17871];
assign MEM[26281] = MEM[14516] + MEM[14915];
assign MEM[26282] = MEM[14518] + MEM[14728];
assign MEM[26283] = MEM[14519] + MEM[14574];
assign MEM[26284] = MEM[14520] + MEM[15599];
assign MEM[26285] = MEM[14521] + MEM[15258];
assign MEM[26286] = MEM[14522] + MEM[15015];
assign MEM[26287] = MEM[14525] + MEM[15852];
assign MEM[26288] = MEM[14527] + MEM[14539];
assign MEM[26289] = MEM[14528] + MEM[14712];
assign MEM[26290] = MEM[14531] + MEM[16963];
assign MEM[26291] = MEM[14533] + MEM[14687];
assign MEM[26292] = MEM[14534] + MEM[16534];
assign MEM[26293] = MEM[14536] + MEM[16026];
assign MEM[26294] = MEM[14537] + MEM[16620];
assign MEM[26295] = MEM[14543] + MEM[18795];
assign MEM[26296] = MEM[14545] + MEM[15028];
assign MEM[26297] = MEM[14547] + MEM[17668];
assign MEM[26298] = MEM[14548] + MEM[17899];
assign MEM[26299] = MEM[14549] + MEM[14851];
assign MEM[26300] = MEM[14550] + MEM[14864];
assign MEM[26301] = MEM[14551] + MEM[15700];
assign MEM[26302] = MEM[14552] + MEM[17439];
assign MEM[26303] = MEM[14553] + MEM[15012];
assign MEM[26304] = MEM[14554] + MEM[18171];
assign MEM[26305] = MEM[14555] + MEM[15672];
assign MEM[26306] = MEM[14557] + MEM[15865];
assign MEM[26307] = MEM[14558] + MEM[18370];
assign MEM[26308] = MEM[14562] + MEM[15510];
assign MEM[26309] = MEM[14563] + MEM[16932];
assign MEM[26310] = MEM[14564] + MEM[16252];
assign MEM[26311] = MEM[14565] + MEM[17501];
assign MEM[26312] = MEM[14566] + MEM[16420];
assign MEM[26313] = MEM[14568] + MEM[16259];
assign MEM[26314] = MEM[14570] + MEM[15087];
assign MEM[26315] = MEM[14571] + MEM[15018];
assign MEM[26316] = MEM[14573] + MEM[16754];
assign MEM[26317] = MEM[14576] + MEM[16955];
assign MEM[26318] = MEM[14578] + MEM[16262];
assign MEM[26319] = MEM[14579] + MEM[16070];
assign MEM[26320] = MEM[14582] + MEM[14839];
assign MEM[26321] = MEM[14590] + MEM[15140];
assign MEM[26322] = MEM[14591] + MEM[15409];
assign MEM[26323] = MEM[14592] + MEM[16035];
assign MEM[26324] = MEM[14593] + MEM[15108];
assign MEM[26325] = MEM[14595] + MEM[15245];
assign MEM[26326] = MEM[14597] + MEM[17416];
assign MEM[26327] = MEM[14598] + MEM[15374];
assign MEM[26328] = MEM[14599] + MEM[14662];
assign MEM[26329] = MEM[14600] + MEM[14651];
assign MEM[26330] = MEM[14603] + MEM[16147];
assign MEM[26331] = MEM[14606] + MEM[14901];
assign MEM[26332] = MEM[14608] + MEM[17720];
assign MEM[26333] = MEM[14609] + MEM[14717];
assign MEM[26334] = MEM[14611] + MEM[16555];
assign MEM[26335] = MEM[14613] + MEM[15788];
assign MEM[26336] = MEM[14615] + MEM[16821];
assign MEM[26337] = MEM[14616] + MEM[17712];
assign MEM[26338] = MEM[14617] + MEM[15827];
assign MEM[26339] = MEM[14618] + MEM[15404];
assign MEM[26340] = MEM[14619] + MEM[17246];
assign MEM[26341] = MEM[14620] + MEM[17356];
assign MEM[26342] = MEM[14624] + MEM[15160];
assign MEM[26343] = MEM[14625] + MEM[20493];
assign MEM[26344] = MEM[14626] + MEM[14922];
assign MEM[26345] = MEM[14627] + MEM[17470];
assign MEM[26346] = MEM[14631] + MEM[15680];
assign MEM[26347] = MEM[14632] + MEM[17017];
assign MEM[26348] = MEM[14633] + MEM[15199];
assign MEM[26349] = MEM[14634] + MEM[15152];
assign MEM[26350] = MEM[14635] + MEM[15860];
assign MEM[26351] = MEM[14637] + MEM[15453];
assign MEM[26352] = MEM[14638] + MEM[16097];
assign MEM[26353] = MEM[14641] + MEM[16957];
assign MEM[26354] = MEM[14644] + MEM[14964];
assign MEM[26355] = MEM[14645] + MEM[16223];
assign MEM[26356] = MEM[14646] + MEM[16280];
assign MEM[26357] = MEM[14647] + MEM[15054];
assign MEM[26358] = MEM[14648] + MEM[15406];
assign MEM[26359] = MEM[14649] + MEM[15440];
assign MEM[26360] = MEM[14650] + MEM[15339];
assign MEM[26361] = MEM[14652] + MEM[14692];
assign MEM[26362] = MEM[14653] + MEM[18580];
assign MEM[26363] = MEM[14654] + MEM[15314];
assign MEM[26364] = MEM[14655] + MEM[14852];
assign MEM[26365] = MEM[14657] + MEM[16425];
assign MEM[26366] = MEM[14661] + MEM[16683];
assign MEM[26367] = MEM[14663] + MEM[17631];
assign MEM[26368] = MEM[14664] + MEM[15405];
assign MEM[26369] = MEM[14665] + MEM[15134];
assign MEM[26370] = MEM[14666] + MEM[17075];
assign MEM[26371] = MEM[14667] + MEM[17382];
assign MEM[26372] = MEM[14668] + MEM[14987];
assign MEM[26373] = MEM[14671] + MEM[17014];
assign MEM[26374] = MEM[14672] + MEM[16514];
assign MEM[26375] = MEM[14673] + MEM[15315];
assign MEM[26376] = MEM[14676] + MEM[14950];
assign MEM[26377] = MEM[14677] + MEM[17773];
assign MEM[26378] = MEM[14678] + MEM[16052];
assign MEM[26379] = MEM[14679] + MEM[16091];
assign MEM[26380] = MEM[14680] + MEM[18833];
assign MEM[26381] = MEM[14682] + MEM[17473];
assign MEM[26382] = MEM[14683] + MEM[17297];
assign MEM[26383] = MEM[14684] + MEM[16242];
assign MEM[26384] = MEM[14686] + MEM[15473];
assign MEM[26385] = MEM[14688] + MEM[16783];
assign MEM[26386] = MEM[14689] + MEM[16169];
assign MEM[26387] = MEM[14690] + MEM[18114];
assign MEM[26388] = MEM[14691] + MEM[14764];
assign MEM[26389] = MEM[14694] + MEM[15249];
assign MEM[26390] = MEM[14696] + MEM[14849];
assign MEM[26391] = MEM[14697] + MEM[17616];
assign MEM[26392] = MEM[14699] + MEM[15627];
assign MEM[26393] = MEM[14700] + MEM[16527];
assign MEM[26394] = MEM[14701] + MEM[15268];
assign MEM[26395] = MEM[14702] + MEM[14733];
assign MEM[26396] = MEM[14703] + MEM[17009];
assign MEM[26397] = MEM[14704] + MEM[17920];
assign MEM[26398] = MEM[14706] + MEM[17970];
assign MEM[26399] = MEM[14707] + MEM[15374];
assign MEM[26400] = MEM[14708] + MEM[15920];
assign MEM[26401] = MEM[14710] + MEM[15193];
assign MEM[26402] = MEM[14711] + MEM[14957];
assign MEM[26403] = MEM[14713] + MEM[16470];
assign MEM[26404] = MEM[14714] + MEM[15452];
assign MEM[26405] = MEM[14715] + MEM[18487];
assign MEM[26406] = MEM[14716] + MEM[16917];
assign MEM[26407] = MEM[14718] + MEM[18998];
assign MEM[26408] = MEM[14720] + MEM[18031];
assign MEM[26409] = MEM[14722] + MEM[17207];
assign MEM[26410] = MEM[14725] + MEM[15664];
assign MEM[26411] = MEM[14726] + MEM[15239];
assign MEM[26412] = MEM[14727] + MEM[18127];
assign MEM[26413] = MEM[14730] + MEM[18886];
assign MEM[26414] = MEM[14732] + MEM[16833];
assign MEM[26415] = MEM[14734] + MEM[17318];
assign MEM[26416] = MEM[14737] + MEM[17330];
assign MEM[26417] = MEM[14740] + MEM[19694];
assign MEM[26418] = MEM[14742] + MEM[16296];
assign MEM[26419] = MEM[14744] + MEM[17313];
assign MEM[26420] = MEM[14745] + MEM[16704];
assign MEM[26421] = MEM[14747] + MEM[16518];
assign MEM[26422] = MEM[14748] + MEM[16595];
assign MEM[26423] = MEM[14751] + MEM[19565];
assign MEM[26424] = MEM[14752] + MEM[14992];
assign MEM[26425] = MEM[14754] + MEM[17181];
assign MEM[26426] = MEM[14756] + MEM[15153];
assign MEM[26427] = MEM[14757] + MEM[15743];
assign MEM[26428] = MEM[14758] + MEM[15103];
assign MEM[26429] = MEM[14760] + MEM[16878];
assign MEM[26430] = MEM[14761] + MEM[16052];
assign MEM[26431] = MEM[14765] + MEM[15221];
assign MEM[26432] = MEM[14766] + MEM[16533];
assign MEM[26433] = MEM[14770] + MEM[15631];
assign MEM[26434] = MEM[14773] + MEM[17422];
assign MEM[26435] = MEM[14774] + MEM[16113];
assign MEM[26436] = MEM[14776] + MEM[19177];
assign MEM[26437] = MEM[14777] + MEM[17966];
assign MEM[26438] = MEM[14778] + MEM[15400];
assign MEM[26439] = MEM[14779] + MEM[17584];
assign MEM[26440] = MEM[14780] + MEM[15788];
assign MEM[26441] = MEM[14782] + MEM[15250];
assign MEM[26442] = MEM[14783] + MEM[16087];
assign MEM[26443] = MEM[14786] + MEM[15033];
assign MEM[26444] = MEM[14787] + MEM[18187];
assign MEM[26445] = MEM[14789] + MEM[17550];
assign MEM[26446] = MEM[14792] + MEM[15780];
assign MEM[26447] = MEM[14795] + MEM[17257];
assign MEM[26448] = MEM[14798] + MEM[16569];
assign MEM[26449] = MEM[14799] + MEM[15925];
assign MEM[26450] = MEM[14801] + MEM[15173];
assign MEM[26451] = MEM[14802] + MEM[16825];
assign MEM[26452] = MEM[14803] + MEM[18480];
assign MEM[26453] = MEM[14805] + MEM[18213];
assign MEM[26454] = MEM[14806] + MEM[14893];
assign MEM[26455] = MEM[14807] + MEM[16504];
assign MEM[26456] = MEM[14810] + MEM[17833];
assign MEM[26457] = MEM[14813] + MEM[17463];
assign MEM[26458] = MEM[14815] + MEM[17649];
assign MEM[26459] = MEM[14816] + MEM[17325];
assign MEM[26460] = MEM[14817] + MEM[14996];
assign MEM[26461] = MEM[14818] + MEM[19512];
assign MEM[26462] = MEM[14821] + MEM[16866];
assign MEM[26463] = MEM[14822] + MEM[15204];
assign MEM[26464] = MEM[14824] + MEM[16223];
assign MEM[26465] = MEM[14825] + MEM[16302];
assign MEM[26466] = MEM[14826] + MEM[15612];
assign MEM[26467] = MEM[14827] + MEM[15895];
assign MEM[26468] = MEM[14828] + MEM[15088];
assign MEM[26469] = MEM[14829] + MEM[15060];
assign MEM[26470] = MEM[14831] + MEM[17924];
assign MEM[26471] = MEM[14833] + MEM[16207];
assign MEM[26472] = MEM[14834] + MEM[17304];
assign MEM[26473] = MEM[14835] + MEM[16277];
assign MEM[26474] = MEM[14836] + MEM[15120];
assign MEM[26475] = MEM[14837] + MEM[20899];
assign MEM[26476] = MEM[14840] + MEM[18234];
assign MEM[26477] = MEM[14841] + MEM[15567];
assign MEM[26478] = MEM[14842] + MEM[16630];
assign MEM[26479] = MEM[14843] + MEM[14935];
assign MEM[26480] = MEM[14846] + MEM[16157];
assign MEM[26481] = MEM[14850] + MEM[18013];
assign MEM[26482] = MEM[14855] + MEM[16389];
assign MEM[26483] = MEM[14856] + MEM[16340];
assign MEM[26484] = MEM[14858] + MEM[16197];
assign MEM[26485] = MEM[14860] + MEM[15784];
assign MEM[26486] = MEM[14861] + MEM[16657];
assign MEM[26487] = MEM[14862] + MEM[17511];
assign MEM[26488] = MEM[14863] + MEM[14903];
assign MEM[26489] = MEM[14866] + MEM[17912];
assign MEM[26490] = MEM[14867] + MEM[16448];
assign MEM[26491] = MEM[14869] + MEM[18522];
assign MEM[26492] = MEM[14872] + MEM[15419];
assign MEM[26493] = MEM[14874] + MEM[17376];
assign MEM[26494] = MEM[14876] + MEM[16289];
assign MEM[26495] = MEM[14878] + MEM[15826];
assign MEM[26496] = MEM[14879] + MEM[15598];
assign MEM[26497] = MEM[14880] + MEM[17382];
assign MEM[26498] = MEM[14883] + MEM[18446];
assign MEM[26499] = MEM[14884] + MEM[18099];
assign MEM[26500] = MEM[14885] + MEM[15127];
assign MEM[26501] = MEM[14886] + MEM[15046];
assign MEM[26502] = MEM[14888] + MEM[17536];
assign MEM[26503] = MEM[14889] + MEM[16632];
assign MEM[26504] = MEM[14892] + MEM[15823];
assign MEM[26505] = MEM[14895] + MEM[15076];
assign MEM[26506] = MEM[14897] + MEM[17549];
assign MEM[26507] = MEM[14905] + MEM[16334];
assign MEM[26508] = MEM[14908] + MEM[16784];
assign MEM[26509] = MEM[14909] + MEM[17619];
assign MEM[26510] = MEM[14910] + MEM[15214];
assign MEM[26511] = MEM[14911] + MEM[15192];
assign MEM[26512] = MEM[14912] + MEM[17521];
assign MEM[26513] = MEM[14914] + MEM[15420];
assign MEM[26514] = MEM[14918] + MEM[16160];
assign MEM[26515] = MEM[14920] + MEM[15426];
assign MEM[26516] = MEM[14921] + MEM[16177];
assign MEM[26517] = MEM[14923] + MEM[16452];
assign MEM[26518] = MEM[14924] + MEM[15078];
assign MEM[26519] = MEM[14925] + MEM[16953];
assign MEM[26520] = MEM[14926] + MEM[15022];
assign MEM[26521] = MEM[14927] + MEM[16818];
assign MEM[26522] = MEM[14928] + MEM[15031];
assign MEM[26523] = MEM[14929] + MEM[17430];
assign MEM[26524] = MEM[14931] + MEM[15645];
assign MEM[26525] = MEM[14934] + MEM[16628];
assign MEM[26526] = MEM[14936] + MEM[19807];
assign MEM[26527] = MEM[14938] + MEM[17502];
assign MEM[26528] = MEM[14939] + MEM[16704];
assign MEM[26529] = MEM[14940] + MEM[15382];
assign MEM[26530] = MEM[14941] + MEM[17515];
assign MEM[26531] = MEM[14943] + MEM[17794];
assign MEM[26532] = MEM[14945] + MEM[15251];
assign MEM[26533] = MEM[14946] + MEM[15318];
assign MEM[26534] = MEM[14947] + MEM[15534];
assign MEM[26535] = MEM[14948] + MEM[15065];
assign MEM[26536] = MEM[14949] + MEM[16228];
assign MEM[26537] = MEM[14953] + MEM[15640];
assign MEM[26538] = MEM[14954] + MEM[17020];
assign MEM[26539] = MEM[14956] + MEM[14995];
assign MEM[26540] = MEM[14958] + MEM[17800];
assign MEM[26541] = MEM[14960] + MEM[18621];
assign MEM[26542] = MEM[14962] + MEM[15196];
assign MEM[26543] = MEM[14963] + MEM[19669];
assign MEM[26544] = MEM[14965] + MEM[16381];
assign MEM[26545] = MEM[14967] + MEM[16078];
assign MEM[26546] = MEM[14968] + MEM[17153];
assign MEM[26547] = MEM[14971] + MEM[17099];
assign MEM[26548] = MEM[14972] + MEM[17569];
assign MEM[26549] = MEM[14973] + MEM[15279];
assign MEM[26550] = MEM[14974] + MEM[16358];
assign MEM[26551] = MEM[14976] + MEM[15444];
assign MEM[26552] = MEM[14978] + MEM[15338];
assign MEM[26553] = MEM[14979] + MEM[14991];
assign MEM[26554] = MEM[14981] + MEM[19827];
assign MEM[26555] = MEM[14982] + MEM[15138];
assign MEM[26556] = MEM[14983] + MEM[16754];
assign MEM[26557] = MEM[14985] + MEM[15267];
assign MEM[26558] = MEM[14993] + MEM[17326];
assign MEM[26559] = MEM[14994] + MEM[15946];
assign MEM[26560] = MEM[14997] + MEM[17947];
assign MEM[26561] = MEM[15001] + MEM[17614];
assign MEM[26562] = MEM[15003] + MEM[16137];
assign MEM[26563] = MEM[15004] + MEM[17143];
assign MEM[26564] = MEM[15005] + MEM[16169];
assign MEM[26565] = MEM[15009] + MEM[17406];
assign MEM[26566] = MEM[15010] + MEM[15066];
assign MEM[26567] = MEM[15013] + MEM[15161];
assign MEM[26568] = MEM[15014] + MEM[17743];
assign MEM[26569] = MEM[15016] + MEM[15212];
assign MEM[26570] = MEM[15019] + MEM[18193];
assign MEM[26571] = MEM[15020] + MEM[16263];
assign MEM[26572] = MEM[15023] + MEM[15384];
assign MEM[26573] = MEM[15026] + MEM[15130];
assign MEM[26574] = MEM[15027] + MEM[16657];
assign MEM[26575] = MEM[15029] + MEM[17761];
assign MEM[26576] = MEM[15030] + MEM[17118];
assign MEM[26577] = MEM[15032] + MEM[15847];
assign MEM[26578] = MEM[15034] + MEM[17442];
assign MEM[26579] = MEM[15035] + MEM[16560];
assign MEM[26580] = MEM[15037] + MEM[16064];
assign MEM[26581] = MEM[15038] + MEM[15416];
assign MEM[26582] = MEM[15039] + MEM[16939];
assign MEM[26583] = MEM[15040] + MEM[16539];
assign MEM[26584] = MEM[15042] + MEM[15435];
assign MEM[26585] = MEM[15045] + MEM[18276];
assign MEM[26586] = MEM[15048] + MEM[16840];
assign MEM[26587] = MEM[15052] + MEM[16588];
assign MEM[26588] = MEM[15055] + MEM[17579];
assign MEM[26589] = MEM[15057] + MEM[17537];
assign MEM[26590] = MEM[15058] + MEM[16535];
assign MEM[26591] = MEM[15059] + MEM[16283];
assign MEM[26592] = MEM[15061] + MEM[18029];
assign MEM[26593] = MEM[15063] + MEM[17745];
assign MEM[26594] = MEM[15068] + MEM[20054];
assign MEM[26595] = MEM[15069] + MEM[16850];
assign MEM[26596] = MEM[15070] + MEM[15133];
assign MEM[26597] = MEM[15071] + MEM[16397];
assign MEM[26598] = MEM[15072] + MEM[16994];
assign MEM[26599] = MEM[15073] + MEM[16809];
assign MEM[26600] = MEM[15075] + MEM[15942];
assign MEM[26601] = MEM[15077] + MEM[16393];
assign MEM[26602] = MEM[15079] + MEM[18406];
assign MEM[26603] = MEM[15082] + MEM[18515];
assign MEM[26604] = MEM[15083] + MEM[16700];
assign MEM[26605] = MEM[15084] + MEM[16750];
assign MEM[26606] = MEM[15086] + MEM[19308];
assign MEM[26607] = MEM[15093] + MEM[15217];
assign MEM[26608] = MEM[15095] + MEM[16028];
assign MEM[26609] = MEM[15099] + MEM[20140];
assign MEM[26610] = MEM[15101] + MEM[16788];
assign MEM[26611] = MEM[15102] + MEM[16188];
assign MEM[26612] = MEM[15104] + MEM[19282];
assign MEM[26613] = MEM[15105] + MEM[18106];
assign MEM[26614] = MEM[15106] + MEM[16786];
assign MEM[26615] = MEM[15109] + MEM[15895];
assign MEM[26616] = MEM[15110] + MEM[15951];
assign MEM[26617] = MEM[15112] + MEM[15520];
assign MEM[26618] = MEM[15113] + MEM[17475];
assign MEM[26619] = MEM[15114] + MEM[16959];
assign MEM[26620] = MEM[15115] + MEM[16095];
assign MEM[26621] = MEM[15118] + MEM[17280];
assign MEM[26622] = MEM[15119] + MEM[16501];
assign MEM[26623] = MEM[15121] + MEM[15261];
assign MEM[26624] = MEM[15122] + MEM[17805];
assign MEM[26625] = MEM[15124] + MEM[16520];
assign MEM[26626] = MEM[15125] + MEM[16078];
assign MEM[26627] = MEM[15128] + MEM[15914];
assign MEM[26628] = MEM[15129] + MEM[17263];
assign MEM[26629] = MEM[15132] + MEM[16296];
assign MEM[26630] = MEM[15135] + MEM[16791];
assign MEM[26631] = MEM[15137] + MEM[15414];
assign MEM[26632] = MEM[15139] + MEM[18040];
assign MEM[26633] = MEM[15142] + MEM[17282];
assign MEM[26634] = MEM[15145] + MEM[16600];
assign MEM[26635] = MEM[15147] + MEM[17296];
assign MEM[26636] = MEM[15148] + MEM[15245];
assign MEM[26637] = MEM[15149] + MEM[18088];
assign MEM[26638] = MEM[15150] + MEM[15202];
assign MEM[26639] = MEM[15155] + MEM[15172];
assign MEM[26640] = MEM[15156] + MEM[16023];
assign MEM[26641] = MEM[15157] + MEM[18177];
assign MEM[26642] = MEM[15158] + MEM[17202];
assign MEM[26643] = MEM[15162] + MEM[18555];
assign MEM[26644] = MEM[15165] + MEM[15746];
assign MEM[26645] = MEM[15168] + MEM[18730];
assign MEM[26646] = MEM[15169] + MEM[17218];
assign MEM[26647] = MEM[15170] + MEM[15801];
assign MEM[26648] = MEM[15175] + MEM[15362];
assign MEM[26649] = MEM[15176] + MEM[15516];
assign MEM[26650] = MEM[15177] + MEM[16846];
assign MEM[26651] = MEM[15178] + MEM[15296];
assign MEM[26652] = MEM[15181] + MEM[15349];
assign MEM[26653] = MEM[15182] + MEM[17988];
assign MEM[26654] = MEM[15185] + MEM[16217];
assign MEM[26655] = MEM[15187] + MEM[19304];
assign MEM[26656] = MEM[15188] + MEM[16450];
assign MEM[26657] = MEM[15189] + MEM[16701];
assign MEM[26658] = MEM[15194] + MEM[16481];
assign MEM[26659] = MEM[15195] + MEM[15276];
assign MEM[26660] = MEM[15197] + MEM[16142];
assign MEM[26661] = MEM[15198] + MEM[16335];
assign MEM[26662] = MEM[15200] + MEM[15717];
assign MEM[26663] = MEM[15205] + MEM[16215];
assign MEM[26664] = MEM[15209] + MEM[15264];
assign MEM[26665] = MEM[15213] + MEM[16571];
assign MEM[26666] = MEM[15215] + MEM[17801];
assign MEM[26667] = MEM[15216] + MEM[19481];
assign MEM[26668] = MEM[15220] + MEM[16587];
assign MEM[26669] = MEM[15222] + MEM[17867];
assign MEM[26670] = MEM[15223] + MEM[16752];
assign MEM[26671] = MEM[15224] + MEM[16640];
assign MEM[26672] = MEM[15225] + MEM[17577];
assign MEM[26673] = MEM[15226] + MEM[17438];
assign MEM[26674] = MEM[15227] + MEM[16759];
assign MEM[26675] = MEM[15229] + MEM[15729];
assign MEM[26676] = MEM[15230] + MEM[15350];
assign MEM[26677] = MEM[15231] + MEM[16878];
assign MEM[26678] = MEM[15232] + MEM[16926];
assign MEM[26679] = MEM[15234] + MEM[18220];
assign MEM[26680] = MEM[15236] + MEM[17339];
assign MEM[26681] = MEM[15238] + MEM[16194];
assign MEM[26682] = MEM[15244] + MEM[17356];
assign MEM[26683] = MEM[15246] + MEM[17687];
assign MEM[26684] = MEM[15247] + MEM[15278];
assign MEM[26685] = MEM[15252] + MEM[16369];
assign MEM[26686] = MEM[15255] + MEM[20539];
assign MEM[26687] = MEM[15256] + MEM[18991];
assign MEM[26688] = MEM[15259] + MEM[18841];
assign MEM[26689] = MEM[15260] + MEM[20366];
assign MEM[26690] = MEM[15263] + MEM[16650];
assign MEM[26691] = MEM[15266] + MEM[15514];
assign MEM[26692] = MEM[15270] + MEM[15776];
assign MEM[26693] = MEM[15271] + MEM[17467];
assign MEM[26694] = MEM[15274] + MEM[15639];
assign MEM[26695] = MEM[15275] + MEM[16703];
assign MEM[26696] = MEM[15277] + MEM[18680];
assign MEM[26697] = MEM[15280] + MEM[17669];
assign MEM[26698] = MEM[15281] + MEM[17683];
assign MEM[26699] = MEM[15282] + MEM[17804];
assign MEM[26700] = MEM[15283] + MEM[18712];
assign MEM[26701] = MEM[15285] + MEM[15366];
assign MEM[26702] = MEM[15287] + MEM[17489];
assign MEM[26703] = MEM[15288] + MEM[15347];
assign MEM[26704] = MEM[15290] + MEM[16809];
assign MEM[26705] = MEM[15291] + MEM[17855];
assign MEM[26706] = MEM[15292] + MEM[15379];
assign MEM[26707] = MEM[15293] + MEM[15313];
assign MEM[26708] = MEM[15294] + MEM[15455];
assign MEM[26709] = MEM[15295] + MEM[16798];
assign MEM[26710] = MEM[15297] + MEM[17442];
assign MEM[26711] = MEM[15302] + MEM[17582];
assign MEM[26712] = MEM[15303] + MEM[17938];
assign MEM[26713] = MEM[15304] + MEM[18379];
assign MEM[26714] = MEM[15305] + MEM[16268];
assign MEM[26715] = MEM[15306] + MEM[17941];
assign MEM[26716] = MEM[15307] + MEM[18426];
assign MEM[26717] = MEM[15308] + MEM[18152];
assign MEM[26718] = MEM[15309] + MEM[15753];
assign MEM[26719] = MEM[15310] + MEM[16542];
assign MEM[26720] = MEM[15312] + MEM[16377];
assign MEM[26721] = MEM[15316] + MEM[16102];
assign MEM[26722] = MEM[15319] + MEM[16892];
assign MEM[26723] = MEM[15320] + MEM[18967];
assign MEM[26724] = MEM[15322] + MEM[16368];
assign MEM[26725] = MEM[15323] + MEM[16632];
assign MEM[26726] = MEM[15324] + MEM[15395];
assign MEM[26727] = MEM[15325] + MEM[16103];
assign MEM[26728] = MEM[15328] + MEM[16438];
assign MEM[26729] = MEM[15329] + MEM[16918];
assign MEM[26730] = MEM[15331] + MEM[15534];
assign MEM[26731] = MEM[15333] + MEM[16840];
assign MEM[26732] = MEM[15334] + MEM[18167];
assign MEM[26733] = MEM[15335] + MEM[16423];
assign MEM[26734] = MEM[15336] + MEM[16813];
assign MEM[26735] = MEM[15337] + MEM[18235];
assign MEM[26736] = MEM[15341] + MEM[17998];
assign MEM[26737] = MEM[15344] + MEM[16577];
assign MEM[26738] = MEM[15345] + MEM[16517];
assign MEM[26739] = MEM[15346] + MEM[17334];
assign MEM[26740] = MEM[15348] + MEM[15750];
assign MEM[26741] = MEM[15352] + MEM[18484];
assign MEM[26742] = MEM[15353] + MEM[16532];
assign MEM[26743] = MEM[15355] + MEM[16196];
assign MEM[26744] = MEM[15357] + MEM[15387];
assign MEM[26745] = MEM[15359] + MEM[16188];
assign MEM[26746] = MEM[15365] + MEM[16764];
assign MEM[26747] = MEM[15367] + MEM[16009];
assign MEM[26748] = MEM[15370] + MEM[16007];
assign MEM[26749] = MEM[15373] + MEM[18066];
assign MEM[26750] = MEM[15376] + MEM[16424];
assign MEM[26751] = MEM[15378] + MEM[16634];
assign MEM[26752] = MEM[15383] + MEM[17146];
assign MEM[26753] = MEM[15388] + MEM[15831];
assign MEM[26754] = MEM[15391] + MEM[17504];
assign MEM[26755] = MEM[15393] + MEM[18888];
assign MEM[26756] = MEM[15394] + MEM[15717];
assign MEM[26757] = MEM[15396] + MEM[15434];
assign MEM[26758] = MEM[15397] + MEM[17092];
assign MEM[26759] = MEM[15398] + MEM[17035];
assign MEM[26760] = MEM[15399] + MEM[17578];
assign MEM[26761] = MEM[15401] + MEM[18397];
assign MEM[26762] = MEM[15410] + MEM[15845];
assign MEM[26763] = MEM[15411] + MEM[17689];
assign MEM[26764] = MEM[15412] + MEM[17067];
assign MEM[26765] = MEM[15413] + MEM[18640];
assign MEM[26766] = MEM[15415] + MEM[17909];
assign MEM[26767] = MEM[15418] + MEM[20378];
assign MEM[26768] = MEM[15421] + MEM[15513];
assign MEM[26769] = MEM[15423] + MEM[16734];
assign MEM[26770] = MEM[15425] + MEM[16142];
assign MEM[26771] = MEM[15428] + MEM[16035];
assign MEM[26772] = MEM[15433] + MEM[15893];
assign MEM[26773] = MEM[15436] + MEM[17507];
assign MEM[26774] = MEM[15443] + MEM[15567];
assign MEM[26775] = MEM[15446] + MEM[17136];
assign MEM[26776] = MEM[15447] + MEM[16427];
assign MEM[26777] = MEM[15448] + MEM[17398];
assign MEM[26778] = MEM[15450] + MEM[16307];
assign MEM[26779] = MEM[15452] + MEM[17072];
assign MEM[26780] = MEM[15453] + MEM[16439];
assign MEM[26781] = MEM[15455] + MEM[16274];
assign MEM[26782] = MEM[15461] + MEM[15723];
assign MEM[26783] = MEM[15471] + MEM[17939];
assign MEM[26784] = MEM[15473] + MEM[18123];
assign MEM[26785] = MEM[15484] + MEM[15813];
assign MEM[26786] = MEM[15489] + MEM[17989];
assign MEM[26787] = MEM[15498] + MEM[16952];
assign MEM[26788] = MEM[15502] + MEM[18536];
assign MEM[26789] = MEM[15503] + MEM[17768];
assign MEM[26790] = MEM[15504] + MEM[18682];
assign MEM[26791] = MEM[15510] + MEM[16891];
assign MEM[26792] = MEM[15514] + MEM[17446];
assign MEM[26793] = MEM[15515] + MEM[16884];
assign MEM[26794] = MEM[15521] + MEM[17777];
assign MEM[26795] = MEM[15531] + MEM[17963];
assign MEM[26796] = MEM[15533] + MEM[16025];
assign MEM[26797] = MEM[15533] + MEM[18602];
assign MEM[26798] = MEM[15535] + MEM[15844];
assign MEM[26799] = MEM[15535] + MEM[17461];
assign MEM[26800] = MEM[15541] + MEM[16481];
assign MEM[26801] = MEM[15541] + MEM[19721];
assign MEM[26802] = MEM[15547] + MEM[17460];
assign MEM[26803] = MEM[15555] + MEM[16285];
assign MEM[26804] = MEM[15562] + MEM[17969];
assign MEM[26805] = MEM[15570] + MEM[17090];
assign MEM[26806] = MEM[15571] + MEM[17402];
assign MEM[26807] = MEM[15572] + MEM[16670];
assign MEM[26808] = MEM[15576] + MEM[16234];
assign MEM[26809] = MEM[15578] + MEM[17651];
assign MEM[26810] = MEM[15591] + MEM[17052];
assign MEM[26811] = MEM[15596] + MEM[16354];
assign MEM[26812] = MEM[15596] + MEM[16456];
assign MEM[26813] = MEM[15599] + MEM[16510];
assign MEM[26814] = MEM[15601] + MEM[16008];
assign MEM[26815] = MEM[15606] + MEM[16603];
assign MEM[26816] = MEM[15607] + MEM[17570];
assign MEM[26817] = MEM[15609] + MEM[17593];
assign MEM[26818] = MEM[15612] + MEM[15860];
assign MEM[26819] = MEM[15617] + MEM[20919];
assign MEM[26820] = MEM[15624] + MEM[17661];
assign MEM[26821] = MEM[15625] + MEM[16436];
assign MEM[26822] = MEM[15631] + MEM[19667];
assign MEM[26823] = MEM[15634] + MEM[16769];
assign MEM[26824] = MEM[15639] + MEM[17523];
assign MEM[26825] = MEM[15646] + MEM[17551];
assign MEM[26826] = MEM[15656] + MEM[16044];
assign MEM[26827] = MEM[15656] + MEM[17575];
assign MEM[26828] = MEM[15660] + MEM[16856];
assign MEM[26829] = MEM[15660] + MEM[17211];
assign MEM[26830] = MEM[15664] + MEM[18046];
assign MEM[26831] = MEM[15665] + MEM[16452];
assign MEM[26832] = MEM[15665] + MEM[18212];
assign MEM[26833] = MEM[15670] + MEM[17857];
assign MEM[26834] = MEM[15672] + MEM[16064];
assign MEM[26835] = MEM[15673] + MEM[16867];
assign MEM[26836] = MEM[15674] + MEM[16731];
assign MEM[26837] = MEM[15680] + MEM[17607];
assign MEM[26838] = MEM[15684] + MEM[15861];
assign MEM[26839] = MEM[15684] + MEM[16575];
assign MEM[26840] = MEM[15689] + MEM[17752];
assign MEM[26841] = MEM[15692] + MEM[16418];
assign MEM[26842] = MEM[15700] + MEM[17737];
assign MEM[26843] = MEM[15702] + MEM[16860];
assign MEM[26844] = MEM[15715] + MEM[17694];
assign MEM[26845] = MEM[15716] + MEM[18456];
assign MEM[26846] = MEM[15723] + MEM[17419];
assign MEM[26847] = MEM[15724] + MEM[17173];
assign MEM[26848] = MEM[15729] + MEM[16439];
assign MEM[26849] = MEM[15743] + MEM[18405];
assign MEM[26850] = MEM[15746] + MEM[17432];
assign MEM[26851] = MEM[15753] + MEM[17176];
assign MEM[26852] = MEM[15756] + MEM[16541];
assign MEM[26853] = MEM[15760] + MEM[16838];
assign MEM[26854] = MEM[15762] + MEM[15826];
assign MEM[26855] = MEM[15770] + MEM[16355];
assign MEM[26856] = MEM[15774] + MEM[16400];
assign MEM[26857] = MEM[15778] + MEM[16788];
assign MEM[26858] = MEM[15778] + MEM[16857];
assign MEM[26859] = MEM[15784] + MEM[16918];
assign MEM[26860] = MEM[15785] + MEM[17663];
assign MEM[26861] = MEM[15787] + MEM[17353];
assign MEM[26862] = MEM[15790] + MEM[16224];
assign MEM[26863] = MEM[15793] + MEM[19608];
assign MEM[26864] = MEM[15801] + MEM[17033];
assign MEM[26865] = MEM[15802] + MEM[16265];
assign MEM[26866] = MEM[15807] + MEM[16685];
assign MEM[26867] = MEM[15808] + MEM[16621];
assign MEM[26868] = MEM[15813] + MEM[16185];
assign MEM[26869] = MEM[15816] + MEM[17063];
assign MEM[26870] = MEM[15819] + MEM[16177];
assign MEM[26871] = MEM[15820] + MEM[19691];
assign MEM[26872] = MEM[15823] + MEM[16157];
assign MEM[26873] = MEM[15827] + MEM[18482];
assign MEM[26874] = MEM[15831] + MEM[17644];
assign MEM[26875] = MEM[15841] + MEM[19029];
assign MEM[26876] = MEM[15847] + MEM[16562];
assign MEM[26877] = MEM[15852] + MEM[16644];
assign MEM[26878] = MEM[15853] + MEM[16402];
assign MEM[26879] = MEM[15865] + MEM[18662];
assign MEM[26880] = MEM[15867] + MEM[17212];
assign MEM[26881] = MEM[15868] + MEM[18070];
assign MEM[26882] = MEM[15871] + MEM[18039];
assign MEM[26883] = MEM[15875] + MEM[19194];
assign MEM[26884] = MEM[15876] + MEM[19297];
assign MEM[26885] = MEM[15886] + MEM[17334];
assign MEM[26886] = MEM[15897] + MEM[18227];
assign MEM[26887] = MEM[15899] + MEM[16538];
assign MEM[26888] = MEM[15903] + MEM[16526];
assign MEM[26889] = MEM[15903] + MEM[17531];
assign MEM[26890] = MEM[15914] + MEM[16733];
assign MEM[26891] = MEM[15920] + MEM[19188];
assign MEM[26892] = MEM[15923] + MEM[17610];
assign MEM[26893] = MEM[15924] + MEM[18051];
assign MEM[26894] = MEM[15925] + MEM[20256];
assign MEM[26895] = MEM[15927] + MEM[17352];
assign MEM[26896] = MEM[15929] + MEM[17647];
assign MEM[26897] = MEM[15931] + MEM[17209];
assign MEM[26898] = MEM[15932] + MEM[17385];
assign MEM[26899] = MEM[15937] + MEM[17780];
assign MEM[26900] = MEM[15938] + MEM[17267];
assign MEM[26901] = MEM[15939] + MEM[17643];
assign MEM[26902] = MEM[15942] + MEM[19138];
assign MEM[26903] = MEM[15946] + MEM[17494];
assign MEM[26904] = MEM[15948] + MEM[19393];
assign MEM[26905] = MEM[15962] + MEM[17950];
assign MEM[26906] = MEM[15963] + MEM[17770];
assign MEM[26907] = MEM[15965] + MEM[17315];
assign MEM[26908] = MEM[15968] + MEM[18575];
assign MEM[26909] = MEM[15974] + MEM[16985];
assign MEM[26910] = MEM[15975] + MEM[17154];
assign MEM[26911] = MEM[15983] + MEM[17513];
assign MEM[26912] = MEM[15984] + MEM[17763];
assign MEM[26913] = MEM[15987] + MEM[16785];
assign MEM[26914] = MEM[15994] + MEM[18140];
assign MEM[26915] = MEM[15995] + MEM[18309];
assign MEM[26916] = MEM[16009] + MEM[17260];
assign MEM[26917] = MEM[16013] + MEM[17496];
assign MEM[26918] = MEM[16018] + MEM[17981];
assign MEM[26919] = MEM[16021] + MEM[16326];
assign MEM[26920] = MEM[16023] + MEM[18931];
assign MEM[26921] = MEM[16026] + MEM[17329];
assign MEM[26922] = MEM[16031] + MEM[16085];
assign MEM[26923] = MEM[16040] + MEM[16767];
assign MEM[26924] = MEM[16044] + MEM[16787];
assign MEM[26925] = MEM[16049] + MEM[18304];
assign MEM[26926] = MEM[16059] + MEM[17851];
assign MEM[26927] = MEM[16061] + MEM[17821];
assign MEM[26928] = MEM[16065] + MEM[18854];
assign MEM[26929] = MEM[16066] + MEM[17403];
assign MEM[26930] = MEM[16070] + MEM[16739];
assign MEM[26931] = MEM[16073] + MEM[16999];
assign MEM[26932] = MEM[16091] + MEM[17862];
assign MEM[26933] = MEM[16094] + MEM[18726];
assign MEM[26934] = MEM[16095] + MEM[18112];
assign MEM[26935] = MEM[16102] + MEM[16962];
assign MEM[26936] = MEM[16103] + MEM[16283];
assign MEM[26937] = MEM[16104] + MEM[17881];
assign MEM[26938] = MEM[16113] + MEM[17958];
assign MEM[26939] = MEM[16117] + MEM[16460];
assign MEM[26940] = MEM[16126] + MEM[19121];
assign MEM[26941] = MEM[16128] + MEM[17173];
assign MEM[26942] = MEM[16128] + MEM[17440];
assign MEM[26943] = MEM[16138] + MEM[17914];
assign MEM[26944] = MEM[16140] + MEM[16266];
assign MEM[26945] = MEM[16140] + MEM[16879];
assign MEM[26946] = MEM[16147] + MEM[16279];
assign MEM[26947] = MEM[16156] + MEM[19617];
assign MEM[26948] = MEM[16160] + MEM[17133];
assign MEM[26949] = MEM[16165] + MEM[16411];
assign MEM[26950] = MEM[16166] + MEM[17908];
assign MEM[26951] = MEM[16171] + MEM[17269];
assign MEM[26952] = MEM[16175] + MEM[18190];
assign MEM[26953] = MEM[16181] + MEM[16954];
assign MEM[26954] = MEM[16183] + MEM[16446];
assign MEM[26955] = MEM[16183] + MEM[17540];
assign MEM[26956] = MEM[16189] + MEM[17038];
assign MEM[26957] = MEM[16190] + MEM[17527];
assign MEM[26958] = MEM[16192] + MEM[16953];
assign MEM[26959] = MEM[16194] + MEM[17673];
assign MEM[26960] = MEM[16195] + MEM[16746];
assign MEM[26961] = MEM[16197] + MEM[16432];
assign MEM[26962] = MEM[16200] + MEM[16968];
assign MEM[26963] = MEM[16203] + MEM[18485];
assign MEM[26964] = MEM[16211] + MEM[16779];
assign MEM[26965] = MEM[16215] + MEM[17171];
assign MEM[26966] = MEM[16217] + MEM[17708];
assign MEM[26967] = MEM[16221] + MEM[17292];
assign MEM[26968] = MEM[16224] + MEM[17954];
assign MEM[26969] = MEM[16233] + MEM[17307];
assign MEM[26970] = MEM[16234] + MEM[17681];
assign MEM[26971] = MEM[16240] + MEM[17354];
assign MEM[26972] = MEM[16242] + MEM[17205];
assign MEM[26973] = MEM[16247] + MEM[18557];
assign MEM[26974] = MEM[16249] + MEM[16694];
assign MEM[26975] = MEM[16249] + MEM[17959];
assign MEM[26976] = MEM[16252] + MEM[17621];
assign MEM[26977] = MEM[16253] + MEM[18887];
assign MEM[26978] = MEM[16255] + MEM[16533];
assign MEM[26979] = MEM[16255] + MEM[16836];
assign MEM[26980] = MEM[16258] + MEM[17990];
assign MEM[26981] = MEM[16259] + MEM[17152];
assign MEM[26982] = MEM[16262] + MEM[19384];
assign MEM[26983] = MEM[16263] + MEM[18567];
assign MEM[26984] = MEM[16265] + MEM[17624];
assign MEM[26985] = MEM[16266] + MEM[17872];
assign MEM[26986] = MEM[16273] + MEM[16366];
assign MEM[26987] = MEM[16274] + MEM[17848];
assign MEM[26988] = MEM[16277] + MEM[20602];
assign MEM[26989] = MEM[16279] + MEM[18977];
assign MEM[26990] = MEM[16280] + MEM[17528];
assign MEM[26991] = MEM[16282] + MEM[17238];
assign MEM[26992] = MEM[16284] + MEM[17113];
assign MEM[26993] = MEM[16285] + MEM[16831];
assign MEM[26994] = MEM[16286] + MEM[20496];
assign MEM[26995] = MEM[16289] + MEM[17815];
assign MEM[26996] = MEM[16293] + MEM[17082];
assign MEM[26997] = MEM[16301] + MEM[17101];
assign MEM[26998] = MEM[16302] + MEM[17338];
assign MEM[26999] = MEM[16307] + MEM[17721];
assign MEM[27000] = MEM[16326] + MEM[16956];
assign MEM[27001] = MEM[16334] + MEM[18165];
assign MEM[27002] = MEM[16335] + MEM[17466];
assign MEM[27003] = MEM[16338] + MEM[17735];
assign MEM[27004] = MEM[16339] + MEM[18085];
assign MEM[27005] = MEM[16340] + MEM[16342];
assign MEM[27006] = MEM[16354] + MEM[18434];
assign MEM[27007] = MEM[16355] + MEM[17819];
assign MEM[27008] = MEM[16358] + MEM[18142];
assign MEM[27009] = MEM[16363] + MEM[17373];
assign MEM[27010] = MEM[16366] + MEM[17239];
assign MEM[27011] = MEM[16367] + MEM[17760];
assign MEM[27012] = MEM[16369] + MEM[17310];
assign MEM[27013] = MEM[16376] + MEM[16778];
assign MEM[27014] = MEM[16376] + MEM[19072];
assign MEM[27015] = MEM[16377] + MEM[17185];
assign MEM[27016] = MEM[16381] + MEM[17829];
assign MEM[27017] = MEM[16388] + MEM[19777];
assign MEM[27018] = MEM[16390] + MEM[17900];
assign MEM[27019] = MEM[16393] + MEM[18579];
assign MEM[27020] = MEM[16394] + MEM[17650];
assign MEM[27021] = MEM[16397] + MEM[18318];
assign MEM[27022] = MEM[16401] + MEM[16499];
assign MEM[27023] = MEM[16403] + MEM[17793];
assign MEM[27024] = MEM[16411] + MEM[17807];
assign MEM[27025] = MEM[16414] + MEM[16927];
assign MEM[27026] = MEM[16414] + MEM[18962];
assign MEM[27027] = MEM[16418] + MEM[17748];
assign MEM[27028] = MEM[16420] + MEM[17547];
assign MEM[27029] = MEM[16423] + MEM[17358];
assign MEM[27030] = MEM[16424] + MEM[19099];
assign MEM[27031] = MEM[16425] + MEM[18274];
assign MEM[27032] = MEM[16427] + MEM[16736];
assign MEM[27033] = MEM[16432] + MEM[19227];
assign MEM[27034] = MEM[16434] + MEM[18472];
assign MEM[27035] = MEM[16436] + MEM[17407];
assign MEM[27036] = MEM[16438] + MEM[19199];
assign MEM[27037] = MEM[16442] + MEM[18008];
assign MEM[27038] = MEM[16446] + MEM[16916];
assign MEM[27039] = MEM[16448] + MEM[16786];
assign MEM[27040] = MEM[16450] + MEM[17991];
assign MEM[27041] = MEM[16456] + MEM[18477];
assign MEM[27042] = MEM[16470] + MEM[17913];
assign MEM[27043] = MEM[16478] + MEM[18868];
assign MEM[27044] = MEM[16484] + MEM[19164];
assign MEM[27045] = MEM[16493] + MEM[17493];
assign MEM[27046] = MEM[16501] + MEM[18157];
assign MEM[27047] = MEM[16502] + MEM[17147];
assign MEM[27048] = MEM[16502] + MEM[17402];
assign MEM[27049] = MEM[16509] + MEM[19080];
assign MEM[27050] = MEM[16510] + MEM[17844];
assign MEM[27051] = MEM[16513] + MEM[16943];
assign MEM[27052] = MEM[16513] + MEM[17636];
assign MEM[27053] = MEM[16514] + MEM[16743];
assign MEM[27054] = MEM[16516] + MEM[18502];
assign MEM[27055] = MEM[16517] + MEM[17266];
assign MEM[27056] = MEM[16520] + MEM[17322];
assign MEM[27057] = MEM[16525] + MEM[20540];
assign MEM[27058] = MEM[16526] + MEM[16573];
assign MEM[27059] = MEM[16527] + MEM[19399];
assign MEM[27060] = MEM[16531] + MEM[17051];
assign MEM[27061] = MEM[16532] + MEM[17222];
assign MEM[27062] = MEM[16534] + MEM[17429];
assign MEM[27063] = MEM[16535] + MEM[18103];
assign MEM[27064] = MEM[16536] + MEM[17273];
assign MEM[27065] = MEM[16539] + MEM[16662];
assign MEM[27066] = MEM[16542] + MEM[23090];
assign MEM[27067] = MEM[16547] + MEM[17447];
assign MEM[27068] = MEM[16548] + MEM[17296];
assign MEM[27069] = MEM[16548] + MEM[19722];
assign MEM[27070] = MEM[16549] + MEM[17378];
assign MEM[27071] = MEM[16549] + MEM[17598];
assign MEM[27072] = MEM[16552] + MEM[18303];
assign MEM[27073] = MEM[16555] + MEM[16790];
assign MEM[27074] = MEM[16560] + MEM[17461];
assign MEM[27075] = MEM[16561] + MEM[17509];
assign MEM[27076] = MEM[16562] + MEM[18353];
assign MEM[27077] = MEM[16563] + MEM[17006];
assign MEM[27078] = MEM[16565] + MEM[17703];
assign MEM[27079] = MEM[16566] + MEM[17102];
assign MEM[27080] = MEM[16566] + MEM[19711];
assign MEM[27081] = MEM[16569] + MEM[17149];
assign MEM[27082] = MEM[16571] + MEM[19214];
assign MEM[27083] = MEM[16573] + MEM[17608];
assign MEM[27084] = MEM[16575] + MEM[18740];
assign MEM[27085] = MEM[16577] + MEM[17751];
assign MEM[27086] = MEM[16579] + MEM[17305];
assign MEM[27087] = MEM[16585] + MEM[18298];
assign MEM[27088] = MEM[16587] + MEM[17524];
assign MEM[27089] = MEM[16588] + MEM[17272];
assign MEM[27090] = MEM[16595] + MEM[17465];
assign MEM[27091] = MEM[16600] + MEM[16914];
assign MEM[27092] = MEM[16602] + MEM[19115];
assign MEM[27093] = MEM[16605] + MEM[16795];
assign MEM[27094] = MEM[16606] + MEM[16636];
assign MEM[27095] = MEM[16606] + MEM[17245];
assign MEM[27096] = MEM[16611] + MEM[16645];
assign MEM[27097] = MEM[16611] + MEM[16846];
assign MEM[27098] = MEM[16612] + MEM[18050];
assign MEM[27099] = MEM[16614] + MEM[17755];
assign MEM[27100] = MEM[16620] + MEM[16932];
assign MEM[27101] = MEM[16621] + MEM[16997];
assign MEM[27102] = MEM[16624] + MEM[19176];
assign MEM[27103] = MEM[16627] + MEM[18811];
assign MEM[27104] = MEM[16628] + MEM[18535];
assign MEM[27105] = MEM[16638] + MEM[16902];
assign MEM[27106] = MEM[16640] + MEM[18067];
assign MEM[27107] = MEM[16644] + MEM[19144];
assign MEM[27108] = MEM[16645] + MEM[17690];
assign MEM[27109] = MEM[16651] + MEM[16935];
assign MEM[27110] = MEM[16651] + MEM[17728];
assign MEM[27111] = MEM[16654] + MEM[17590];
assign MEM[27112] = MEM[16654] + MEM[17698];
assign MEM[27113] = MEM[16656] + MEM[18291];
assign MEM[27114] = MEM[16662] + MEM[18620];
assign MEM[27115] = MEM[16665] + MEM[17061];
assign MEM[27116] = MEM[16665] + MEM[17411];
assign MEM[27117] = MEM[16670] + MEM[16831];
assign MEM[27118] = MEM[16683] + MEM[17150];
assign MEM[27119] = MEM[16685] + MEM[17674];
assign MEM[27120] = MEM[16686] + MEM[17202];
assign MEM[27121] = MEM[16691] + MEM[17823];
assign MEM[27122] = MEM[16694] + MEM[20235];
assign MEM[27123] = MEM[16695] + MEM[17790];
assign MEM[27124] = MEM[16700] + MEM[19754];
assign MEM[27125] = MEM[16702] + MEM[17423];
assign MEM[27126] = MEM[16703] + MEM[18181];
assign MEM[27127] = MEM[16711] + MEM[18175];
assign MEM[27128] = MEM[16718] + MEM[16864];
assign MEM[27129] = MEM[16718] + MEM[18802];
assign MEM[27130] = MEM[16723] + MEM[17542];
assign MEM[27131] = MEM[16731] + MEM[17831];
assign MEM[27132] = MEM[16734] + MEM[19911];
assign MEM[27133] = MEM[16736] + MEM[18153];
assign MEM[27134] = MEM[16738] + MEM[17121];
assign MEM[27135] = MEM[16739] + MEM[18930];
assign MEM[27136] = MEM[16740] + MEM[18464];
assign MEM[27137] = MEM[16741] + MEM[18745];
assign MEM[27138] = MEM[16743] + MEM[18251];
assign MEM[27139] = MEM[16746] + MEM[17830];
assign MEM[27140] = MEM[16750] + MEM[16967];
assign MEM[27141] = MEM[16752] + MEM[19266];
assign MEM[27142] = MEM[16762] + MEM[17041];
assign MEM[27143] = MEM[16767] + MEM[17785];
assign MEM[27144] = MEM[16768] + MEM[17046];
assign MEM[27145] = MEM[16768] + MEM[17115];
assign MEM[27146] = MEM[16769] + MEM[19713];
assign MEM[27147] = MEM[16777] + MEM[18608];
assign MEM[27148] = MEM[16778] + MEM[18245];
assign MEM[27149] = MEM[16780] + MEM[17203];
assign MEM[27150] = MEM[16780] + MEM[18481];
assign MEM[27151] = MEM[16783] + MEM[21836];
assign MEM[27152] = MEM[16784] + MEM[17227];
assign MEM[27153] = MEM[16785] + MEM[17149];
assign MEM[27154] = MEM[16787] + MEM[18059];
assign MEM[27155] = MEM[16791] + MEM[17711];
assign MEM[27156] = MEM[16795] + MEM[17533];
assign MEM[27157] = MEM[16796] + MEM[18208];
assign MEM[27158] = MEM[16798] + MEM[17847];
assign MEM[27159] = MEM[16813] + MEM[17075];
assign MEM[27160] = MEM[16818] + MEM[18093];
assign MEM[27161] = MEM[16821] + MEM[18374];
assign MEM[27162] = MEM[16823] + MEM[17736];
assign MEM[27163] = MEM[16823] + MEM[17854];
assign MEM[27164] = MEM[16825] + MEM[17052];
assign MEM[27165] = MEM[16833] + MEM[17982];
assign MEM[27166] = MEM[16836] + MEM[18117];
assign MEM[27167] = MEM[16838] + MEM[17353];
assign MEM[27168] = MEM[16839] + MEM[17445];
assign MEM[27169] = MEM[16839] + MEM[19381];
assign MEM[27170] = MEM[16847] + MEM[17679];
assign MEM[27171] = MEM[16848] + MEM[16963];
assign MEM[27172] = MEM[16848] + MEM[17727];
assign MEM[27173] = MEM[16850] + MEM[19015];
assign MEM[27174] = MEM[16856] + MEM[17227];
assign MEM[27175] = MEM[16857] + MEM[17592];
assign MEM[27176] = MEM[16860] + MEM[17500];
assign MEM[27177] = MEM[16865] + MEM[18305];
assign MEM[27178] = MEM[16866] + MEM[17940];
assign MEM[27179] = MEM[16868] + MEM[17041];
assign MEM[27180] = MEM[16872] + MEM[17765];
assign MEM[27181] = MEM[16879] + MEM[17571];
assign MEM[27182] = MEM[16884] + MEM[17739];
assign MEM[27183] = MEM[16891] + MEM[18976];
assign MEM[27184] = MEM[16892] + MEM[19019];
assign MEM[27185] = MEM[16894] + MEM[17365];
assign MEM[27186] = MEM[16894] + MEM[17517];
assign MEM[27187] = MEM[16902] + MEM[18100];
assign MEM[27188] = MEM[16908] + MEM[20145];
assign MEM[27189] = MEM[16911] + MEM[18691];
assign MEM[27190] = MEM[16912] + MEM[17994];
assign MEM[27191] = MEM[16915] + MEM[17486];
assign MEM[27192] = MEM[16916] + MEM[18789];
assign MEM[27193] = MEM[16917] + MEM[17879];
assign MEM[27194] = MEM[16927] + MEM[17942];
assign MEM[27195] = MEM[16935] + MEM[17470];
assign MEM[27196] = MEM[16939] + MEM[19200];
assign MEM[27197] = MEM[16943] + MEM[17104];
assign MEM[27198] = MEM[16952] + MEM[18164];
assign MEM[27199] = MEM[16955] + MEM[18398];
assign MEM[27200] = MEM[16956] + MEM[19076];
assign MEM[27201] = MEM[16957] + MEM[18445];
assign MEM[27202] = MEM[16958] + MEM[18247];
assign MEM[27203] = MEM[16959] + MEM[17398];
assign MEM[27204] = MEM[16961] + MEM[17427];
assign MEM[27205] = MEM[16962] + MEM[17465];
assign MEM[27206] = MEM[16967] + MEM[17205];
assign MEM[27207] = MEM[16968] + MEM[18236];
assign MEM[27208] = MEM[16985] + MEM[18523];
assign MEM[27209] = MEM[16987] + MEM[17304];
assign MEM[27210] = MEM[16989] + MEM[17818];
assign MEM[27211] = MEM[16994] + MEM[20914];
assign MEM[27212] = MEM[16996] + MEM[17290];
assign MEM[27213] = MEM[16996] + MEM[17652];
assign MEM[27214] = MEM[16999] + MEM[20477];
assign MEM[27215] = MEM[17002] + MEM[17323];
assign MEM[27216] = MEM[17002] + MEM[17634];
assign MEM[27217] = MEM[17006] + MEM[18945];
assign MEM[27218] = MEM[17007] + MEM[18919];
assign MEM[27219] = MEM[17009] + MEM[17123];
assign MEM[27220] = MEM[17013] + MEM[21232];
assign MEM[27221] = MEM[17014] + MEM[18458];
assign MEM[27222] = MEM[17019] + MEM[17029];
assign MEM[27223] = MEM[17020] + MEM[17601];
assign MEM[27224] = MEM[17024] + MEM[17404];
assign MEM[27225] = MEM[17028] + MEM[17568];
assign MEM[27226] = MEM[17028] + MEM[20757];
assign MEM[27227] = MEM[17032] + MEM[17779];
assign MEM[27228] = MEM[17033] + MEM[17480];
assign MEM[27229] = MEM[17035] + MEM[17635];
assign MEM[27230] = MEM[17038] + MEM[18256];
assign MEM[27231] = MEM[17045] + MEM[19083];
assign MEM[27232] = MEM[17046] + MEM[18170];
assign MEM[27233] = MEM[17050] + MEM[18058];
assign MEM[27234] = MEM[17053] + MEM[17401];
assign MEM[27235] = MEM[17054] + MEM[17993];
assign MEM[27236] = MEM[17056] + MEM[17308];
assign MEM[27237] = MEM[17058] + MEM[19891];
assign MEM[27238] = MEM[17061] + MEM[21114];
assign MEM[27239] = MEM[17063] + MEM[18537];
assign MEM[27240] = MEM[17065] + MEM[17452];
assign MEM[27241] = MEM[17067] + MEM[17358];
assign MEM[27242] = MEM[17068] + MEM[17597];
assign MEM[27243] = MEM[17068] + MEM[17895];
assign MEM[27244] = MEM[17072] + MEM[18706];
assign MEM[27245] = MEM[17083] + MEM[17491];
assign MEM[27246] = MEM[17083] + MEM[17820];
assign MEM[27247] = MEM[17084] + MEM[17387];
assign MEM[27248] = MEM[17084] + MEM[20462];
assign MEM[27249] = MEM[17085] + MEM[17463];
assign MEM[27250] = MEM[17085] + MEM[18362];
assign MEM[27251] = MEM[17090] + MEM[19800];
assign MEM[27252] = MEM[17092] + MEM[18323];
assign MEM[27253] = MEM[17093] + MEM[18732];
assign MEM[27254] = MEM[17097] + MEM[18095];
assign MEM[27255] = MEM[17097] + MEM[18603];
assign MEM[27256] = MEM[17099] + MEM[18041];
assign MEM[27257] = MEM[17101] + MEM[18018];
assign MEM[27258] = MEM[17102] + MEM[18817];
assign MEM[27259] = MEM[17113] + MEM[17612];
assign MEM[27260] = MEM[17115] + MEM[20944];
assign MEM[27261] = MEM[17118] + MEM[19765];
assign MEM[27262] = MEM[17121] + MEM[17368];
assign MEM[27263] = MEM[17122] + MEM[17328];
assign MEM[27264] = MEM[17123] + MEM[17928];
assign MEM[27265] = MEM[17125] + MEM[18604];
assign MEM[27266] = MEM[17133] + MEM[17953];
assign MEM[27267] = MEM[17134] + MEM[17146];
assign MEM[27268] = MEM[17134] + MEM[18717];
assign MEM[27269] = MEM[17143] + MEM[18080];
assign MEM[27270] = MEM[17147] + MEM[19137];
assign MEM[27271] = MEM[17150] + MEM[17376];
assign MEM[27272] = MEM[17152] + MEM[19997];
assign MEM[27273] = MEM[17153] + MEM[19720];
assign MEM[27274] = MEM[17154] + MEM[17319];
assign MEM[27275] = MEM[17169] + MEM[17312];
assign MEM[27276] = MEM[17169] + MEM[18194];
assign MEM[27277] = MEM[17170] + MEM[17841];
assign MEM[27278] = MEM[17171] + MEM[18916];
assign MEM[27279] = MEM[17176] + MEM[17659];
assign MEM[27280] = MEM[17179] + MEM[17692];
assign MEM[27281] = MEM[17179] + MEM[18615];
assign MEM[27282] = MEM[17180] + MEM[18875];
assign MEM[27283] = MEM[17181] + MEM[21543];
assign MEM[27284] = MEM[17190] + MEM[18009];
assign MEM[27285] = MEM[17197] + MEM[18573];
assign MEM[27286] = MEM[17198] + MEM[17664];
assign MEM[27287] = MEM[17200] + MEM[17434];
assign MEM[27288] = MEM[17200] + MEM[18520];
assign MEM[27289] = MEM[17201] + MEM[18054];
assign MEM[27290] = MEM[17203] + MEM[17858];
assign MEM[27291] = MEM[17207] + MEM[17333];
assign MEM[27292] = MEM[17209] + MEM[17211];
assign MEM[27293] = MEM[17212] + MEM[17580];
assign MEM[27294] = MEM[17214] + MEM[17685];
assign MEM[27295] = MEM[17214] + MEM[18663];
assign MEM[27296] = MEM[17222] + MEM[17873];
assign MEM[27297] = MEM[17237] + MEM[19501];
assign MEM[27298] = MEM[17238] + MEM[17613];
assign MEM[27299] = MEM[17239] + MEM[17753];
assign MEM[27300] = MEM[17245] + MEM[18373];
assign MEM[27301] = MEM[17246] + MEM[18766];
assign MEM[27302] = MEM[17257] + MEM[18879];
assign MEM[27303] = MEM[17260] + MEM[20988];
assign MEM[27304] = MEM[17262] + MEM[18130];
assign MEM[27305] = MEM[17263] + MEM[22344];
assign MEM[27306] = MEM[17264] + MEM[17436];
assign MEM[27307] = MEM[17264] + MEM[17733];
assign MEM[27308] = MEM[17266] + MEM[18252];
assign MEM[27309] = MEM[17267] + MEM[17587];
assign MEM[27310] = MEM[17269] + MEM[18168];
assign MEM[27311] = MEM[17272] + MEM[17836];
assign MEM[27312] = MEM[17280] + MEM[17791];
assign MEM[27313] = MEM[17282] + MEM[17365];
assign MEM[27314] = MEM[17284] + MEM[18205];
assign MEM[27315] = MEM[17286] + MEM[18533];
assign MEM[27316] = MEM[17292] + MEM[20564];
assign MEM[27317] = MEM[17297] + MEM[17332];
assign MEM[27318] = MEM[17298] + MEM[18401];
assign MEM[27319] = MEM[17305] + MEM[17475];
assign MEM[27320] = MEM[17307] + MEM[18083];
assign MEM[27321] = MEM[17308] + MEM[20821];
assign MEM[27322] = MEM[17310] + MEM[18491];
assign MEM[27323] = MEM[17312] + MEM[18321];
assign MEM[27324] = MEM[17313] + MEM[18561];
assign MEM[27325] = MEM[17315] + MEM[18010];
assign MEM[27326] = MEM[17318] + MEM[19419];
assign MEM[27327] = MEM[17319] + MEM[18364];
assign MEM[27328] = MEM[17322] + MEM[17626];
assign MEM[27329] = MEM[17323] + MEM[17896];
assign MEM[27330] = MEM[17325] + MEM[18134];
assign MEM[27331] = MEM[17328] + MEM[18022];
assign MEM[27332] = MEM[17329] + MEM[18501];
assign MEM[27333] = MEM[17330] + MEM[18935];
assign MEM[27334] = MEM[17332] + MEM[19085];
assign MEM[27335] = MEM[17333] + MEM[17383];
assign MEM[27336] = MEM[17338] + MEM[17766];
assign MEM[27337] = MEM[17339] + MEM[19159];
assign MEM[27338] = MEM[17349] + MEM[18217];
assign MEM[27339] = MEM[17349] + MEM[18729];
assign MEM[27340] = MEM[17352] + MEM[18075];
assign MEM[27341] = MEM[17354] + MEM[18655];
assign MEM[27342] = MEM[17364] + MEM[18437];
assign MEM[27343] = MEM[17368] + MEM[18286];
assign MEM[27344] = MEM[17369] + MEM[17503];
assign MEM[27345] = MEM[17369] + MEM[17925];
assign MEM[27346] = MEM[17370] + MEM[18915];
assign MEM[27347] = MEM[17373] + MEM[17901];
assign MEM[27348] = MEM[17378] + MEM[17922];
assign MEM[27349] = MEM[17379] + MEM[17424];
assign MEM[27350] = MEM[17379] + MEM[17987];
assign MEM[27351] = MEM[17385] + MEM[18347];
assign MEM[27352] = MEM[17387] + MEM[18652];
assign MEM[27353] = MEM[17403] + MEM[18440];
assign MEM[27354] = MEM[17404] + MEM[19710];
assign MEM[27355] = MEM[17405] + MEM[17595];
assign MEM[27356] = MEM[17405] + MEM[18355];
assign MEM[27357] = MEM[17406] + MEM[18566];
assign MEM[27358] = MEM[17407] + MEM[18378];
assign MEM[27359] = MEM[17411] + MEM[17648];
assign MEM[27360] = MEM[17412] + MEM[17428];
assign MEM[27361] = MEM[17412] + MEM[18159];
assign MEM[27362] = MEM[17416] + MEM[19618];
assign MEM[27363] = MEM[17417] + MEM[17572];
assign MEM[27364] = MEM[17417] + MEM[19295];
assign MEM[27365] = MEM[17419] + MEM[19491];
assign MEM[27366] = MEM[17424] + MEM[17825];
assign MEM[27367] = MEM[17430] + MEM[18030];
assign MEM[27368] = MEM[17432] + MEM[19165];
assign MEM[27369] = MEM[17434] + MEM[18173];
assign MEM[27370] = MEM[17436] + MEM[18284];
assign MEM[27371] = MEM[17438] + MEM[18733];
assign MEM[27372] = MEM[17439] + MEM[18238];
assign MEM[27373] = MEM[17440] + MEM[19376];
assign MEM[27374] = MEM[17441] + MEM[17658];
assign MEM[27375] = MEM[17441] + MEM[20052];
assign MEM[27376] = MEM[17445] + MEM[18136];
assign MEM[27377] = MEM[17446] + MEM[17555];
assign MEM[27378] = MEM[17447] + MEM[18693];
assign MEM[27379] = MEM[17452] + MEM[17882];
assign MEM[27380] = MEM[17456] + MEM[17557];
assign MEM[27381] = MEM[17456] + MEM[18722];
assign MEM[27382] = MEM[17460] + MEM[18596];
assign MEM[27383] = MEM[17466] + MEM[18684];
assign MEM[27384] = MEM[17467] + MEM[20479];
assign MEM[27385] = MEM[17474] + MEM[19101];
assign MEM[27386] = MEM[17479] + MEM[18061];
assign MEM[27387] = MEM[17481] + MEM[17849];
assign MEM[27388] = MEM[17484] + MEM[17774];
assign MEM[27389] = MEM[17487] + MEM[17581];
assign MEM[27390] = MEM[17490] + MEM[17722];
assign MEM[27391] = MEM[17492] + MEM[17957];
assign MEM[27392] = MEM[17495] + MEM[18037];
assign MEM[27393] = MEM[17497] + MEM[18063];
assign MEM[27394] = MEM[17499] + MEM[19317];
assign MEM[27395] = MEM[17505] + MEM[18694];
assign MEM[27396] = MEM[17508] + MEM[17814];
assign MEM[27397] = MEM[17514] + MEM[17530];
assign MEM[27398] = MEM[17516] + MEM[17656];
assign MEM[27399] = MEM[17520] + MEM[18182];
assign MEM[27400] = MEM[17522] + MEM[17918];
assign MEM[27401] = MEM[17525] + MEM[18271];
assign MEM[27402] = MEM[17538] + MEM[17926];
assign MEM[27403] = MEM[17541] + MEM[17834];
assign MEM[27404] = MEM[17543] + MEM[18660];
assign MEM[27405] = MEM[17544] + MEM[17824];
assign MEM[27406] = MEM[17545] + MEM[17546];
assign MEM[27407] = MEM[17548] + MEM[17828];
assign MEM[27408] = MEM[17553] + MEM[17628];
assign MEM[27409] = MEM[17560] + MEM[17657];
assign MEM[27410] = MEM[17562] + MEM[17845];
assign MEM[27411] = MEM[17564] + MEM[19096];
assign MEM[27412] = MEM[17574] + MEM[17802];
assign MEM[27413] = MEM[17583] + MEM[18144];
assign MEM[27414] = MEM[17586] + MEM[18606];
assign MEM[27415] = MEM[17589] + MEM[18098];
assign MEM[27416] = MEM[17591] + MEM[17890];
assign MEM[27417] = MEM[17594] + MEM[18311];
assign MEM[27418] = MEM[17599] + MEM[17898];
assign MEM[27419] = MEM[17603] + MEM[17706];
assign MEM[27420] = MEM[17604] + MEM[17654];
assign MEM[27421] = MEM[17605] + MEM[17622];
assign MEM[27422] = MEM[17606] + MEM[17617];
assign MEM[27423] = MEM[17609] + MEM[17700];
assign MEM[27424] = MEM[17611] + MEM[18385];
assign MEM[27425] = MEM[17630] + MEM[17640];
assign MEM[27426] = MEM[17633] + MEM[18087];
assign MEM[27427] = MEM[17637] + MEM[17784];
assign MEM[27428] = MEM[17638] + MEM[17677];
assign MEM[27429] = MEM[17655] + MEM[18433];
assign MEM[27430] = MEM[17660] + MEM[17892];
assign MEM[27431] = MEM[17665] + MEM[17789];
assign MEM[27432] = MEM[17670] + MEM[18320];
assign MEM[27433] = MEM[17671] + MEM[17875];
assign MEM[27434] = MEM[17678] + MEM[18275];
assign MEM[27435] = MEM[17680] + MEM[18264];
assign MEM[27436] = MEM[17682] + MEM[18431];
assign MEM[27437] = MEM[17684] + MEM[17719];
assign MEM[27438] = MEM[17686] + MEM[17726];
assign MEM[27439] = MEM[17691] + MEM[17838];
assign MEM[27440] = MEM[17697] + MEM[18332];
assign MEM[27441] = MEM[17701] + MEM[18176];
assign MEM[27442] = MEM[17704] + MEM[17729];
assign MEM[27443] = MEM[17714] + MEM[18068];
assign MEM[27444] = MEM[17715] + MEM[18005];
assign MEM[27445] = MEM[17717] + MEM[17916];
assign MEM[27446] = MEM[17718] + MEM[18852];
assign MEM[27447] = MEM[17724] + MEM[17952];
assign MEM[27448] = MEM[17741] + MEM[17781];
assign MEM[27449] = MEM[17744] + MEM[18570];
assign MEM[27450] = MEM[17746] + MEM[17972];
assign MEM[27451] = MEM[17749] + MEM[18308];
assign MEM[27452] = MEM[17762] + MEM[18101];
assign MEM[27453] = MEM[17764] + MEM[17856];
assign MEM[27454] = MEM[17767] + MEM[18384];
assign MEM[27455] = MEM[17771] + MEM[17961];
assign MEM[27456] = MEM[17772] + MEM[17843];
assign MEM[27457] = MEM[17775] + MEM[18065];
assign MEM[27458] = MEM[17776] + MEM[17984];
assign MEM[27459] = MEM[17783] + MEM[18721];
assign MEM[27460] = MEM[17787] + MEM[18129];
assign MEM[27461] = MEM[17788] + MEM[17944];
assign MEM[27462] = MEM[17792] + MEM[17889];
assign MEM[27463] = MEM[17795] + MEM[17919];
assign MEM[27464] = MEM[17797] + MEM[18813];
assign MEM[27465] = MEM[17798] + MEM[18390];
assign MEM[27466] = MEM[17803] + MEM[18138];
assign MEM[27467] = MEM[17809] + MEM[18126];
assign MEM[27468] = MEM[17810] + MEM[19134];
assign MEM[27469] = MEM[17811] + MEM[18133];
assign MEM[27470] = MEM[17817] + MEM[18269];
assign MEM[27471] = MEM[17835] + MEM[17978];
assign MEM[27472] = MEM[17837] + MEM[18342];
assign MEM[27473] = MEM[17840] + MEM[18871];
assign MEM[27474] = MEM[17846] + MEM[18735];
assign MEM[27475] = MEM[17859] + MEM[17974];
assign MEM[27476] = MEM[17860] + MEM[17863];
assign MEM[27477] = MEM[17869] + MEM[18294];
assign MEM[27478] = MEM[17870] + MEM[18516];
assign MEM[27479] = MEM[17874] + MEM[18359];
assign MEM[27480] = MEM[17876] + MEM[18563];
assign MEM[27481] = MEM[17878] + MEM[18435];
assign MEM[27482] = MEM[17880] + MEM[18556];
assign MEM[27483] = MEM[17883] + MEM[18178];
assign MEM[27484] = MEM[17885] + MEM[18214];
assign MEM[27485] = MEM[17887] + MEM[18622];
assign MEM[27486] = MEM[17891] + MEM[18279];
assign MEM[27487] = MEM[17893] + MEM[18777];
assign MEM[27488] = MEM[17904] + MEM[18216];
assign MEM[27489] = MEM[17906] + MEM[18016];
assign MEM[27490] = MEM[17910] + MEM[18979];
assign MEM[27491] = MEM[17915] + MEM[18300];
assign MEM[27492] = MEM[17927] + MEM[17971];
assign MEM[27493] = MEM[17929] + MEM[18643];
assign MEM[27494] = MEM[17931] + MEM[18042];
assign MEM[27495] = MEM[17932] + MEM[18237];
assign MEM[27496] = MEM[17933] + MEM[18113];
assign MEM[27497] = MEM[17936] + MEM[18141];
assign MEM[27498] = MEM[17946] + MEM[18012];
assign MEM[27499] = MEM[17948] + MEM[18250];
assign MEM[27500] = MEM[17949] + MEM[18086];
assign MEM[27501] = MEM[17951] + MEM[18062];
assign MEM[27502] = MEM[17955] + MEM[17968];
assign MEM[27503] = MEM[17960] + MEM[18490];
assign MEM[27504] = MEM[17962] + MEM[18226];
assign MEM[27505] = MEM[17964] + MEM[18329];
assign MEM[27506] = MEM[17965] + MEM[18774];
assign MEM[27507] = MEM[17967] + MEM[18702];
assign MEM[27508] = MEM[17975] + MEM[18000];
assign MEM[27509] = MEM[17980] + MEM[18785];
assign MEM[27510] = MEM[17983] + MEM[18121];
assign MEM[27511] = MEM[17985] + MEM[18549];
assign MEM[27512] = MEM[17986] + MEM[18576];
assign MEM[27513] = MEM[17995] + MEM[18736];
assign MEM[27514] = MEM[17997] + MEM[18872];
assign MEM[27515] = MEM[17999] + MEM[18262];
assign MEM[27516] = MEM[18001] + MEM[18191];
assign MEM[27517] = MEM[18003] + MEM[18259];
assign MEM[27518] = MEM[18006] + MEM[18494];
assign MEM[27519] = MEM[18011] + MEM[18407];
assign MEM[27520] = MEM[18014] + MEM[18221];
assign MEM[27521] = MEM[18015] + MEM[18233];
assign MEM[27522] = MEM[18019] + MEM[18218];
assign MEM[27523] = MEM[18021] + MEM[18097];
assign MEM[27524] = MEM[18023] + MEM[20008];
assign MEM[27525] = MEM[18024] + MEM[20342];
assign MEM[27526] = MEM[18025] + MEM[18033];
assign MEM[27527] = MEM[18026] + MEM[18203];
assign MEM[27528] = MEM[18027] + MEM[19009];
assign MEM[27529] = MEM[18032] + MEM[18072];
assign MEM[27530] = MEM[18034] + MEM[18202];
assign MEM[27531] = MEM[18035] + MEM[18757];
assign MEM[27532] = MEM[18036] + MEM[18199];
assign MEM[27533] = MEM[18038] + MEM[18896];
assign MEM[27534] = MEM[18044] + MEM[18400];
assign MEM[27535] = MEM[18045] + MEM[18350];
assign MEM[27536] = MEM[18048] + MEM[19556];
assign MEM[27537] = MEM[18052] + MEM[18334];
assign MEM[27538] = MEM[18053] + MEM[18091];
assign MEM[27539] = MEM[18056] + MEM[18224];
assign MEM[27540] = MEM[18057] + MEM[18442];
assign MEM[27541] = MEM[18060] + MEM[18424];
assign MEM[27542] = MEM[18064] + MEM[18999];
assign MEM[27543] = MEM[18071] + MEM[18780];
assign MEM[27544] = MEM[18074] + MEM[18244];
assign MEM[27545] = MEM[18077] + MEM[18301];
assign MEM[27546] = MEM[18078] + MEM[18387];
assign MEM[27547] = MEM[18084] + MEM[18679];
assign MEM[27548] = MEM[18090] + MEM[18180];
assign MEM[27549] = MEM[18092] + MEM[18287];
assign MEM[27550] = MEM[18105] + MEM[18369];
assign MEM[27551] = MEM[18107] + MEM[18375];
assign MEM[27552] = MEM[18110] + MEM[18568];
assign MEM[27553] = MEM[18111] + MEM[18312];
assign MEM[27554] = MEM[18115] + MEM[18452];
assign MEM[27555] = MEM[18118] + MEM[18461];
assign MEM[27556] = MEM[18125] + MEM[18278];
assign MEM[27557] = MEM[18128] + MEM[18314];
assign MEM[27558] = MEM[18131] + MEM[18357];
assign MEM[27559] = MEM[18135] + MEM[18463];
assign MEM[27560] = MEM[18137] + MEM[18741];
assign MEM[27561] = MEM[18145] + MEM[18667];
assign MEM[27562] = MEM[18146] + MEM[18249];
assign MEM[27563] = MEM[18149] + MEM[19127];
assign MEM[27564] = MEM[18150] + MEM[18209];
assign MEM[27565] = MEM[18154] + MEM[18222];
assign MEM[27566] = MEM[18156] + MEM[19521];
assign MEM[27567] = MEM[18160] + MEM[18169];
assign MEM[27568] = MEM[18161] + MEM[19759];
assign MEM[27569] = MEM[18162] + MEM[18913];
assign MEM[27570] = MEM[18163] + MEM[18189];
assign MEM[27571] = MEM[18172] + MEM[18467];
assign MEM[27572] = MEM[18179] + MEM[18451];
assign MEM[27573] = MEM[18186] + MEM[18995];
assign MEM[27574] = MEM[18188] + MEM[19434];
assign MEM[27575] = MEM[18192] + MEM[18842];
assign MEM[27576] = MEM[18196] + MEM[18688];
assign MEM[27577] = MEM[18197] + MEM[18518];
assign MEM[27578] = MEM[18198] + MEM[18299];
assign MEM[27579] = MEM[18200] + MEM[18246];
assign MEM[27580] = MEM[18201] + MEM[18345];
assign MEM[27581] = MEM[18204] + MEM[18992];
assign MEM[27582] = MEM[18206] + MEM[18917];
assign MEM[27583] = MEM[18207] + MEM[18946];
assign MEM[27584] = MEM[18211] + MEM[18239];
assign MEM[27585] = MEM[18215] + MEM[18302];
assign MEM[27586] = MEM[18219] + MEM[18263];
assign MEM[27587] = MEM[18225] + MEM[18402];
assign MEM[27588] = MEM[18229] + MEM[18687];
assign MEM[27589] = MEM[18230] + MEM[18856];
assign MEM[27590] = MEM[18232] + MEM[18587];
assign MEM[27591] = MEM[18242] + MEM[18619];
assign MEM[27592] = MEM[18248] + MEM[18532];
assign MEM[27593] = MEM[18253] + MEM[18552];
assign MEM[27594] = MEM[18257] + MEM[18657];
assign MEM[27595] = MEM[18266] + MEM[18478];
assign MEM[27596] = MEM[18267] + MEM[18360];
assign MEM[27597] = MEM[18268] + MEM[18755];
assign MEM[27598] = MEM[18270] + MEM[18343];
assign MEM[27599] = MEM[18272] + MEM[18961];
assign MEM[27600] = MEM[18273] + MEM[18819];
assign MEM[27601] = MEM[18277] + MEM[18763];
assign MEM[27602] = MEM[18280] + MEM[19203];
assign MEM[27603] = MEM[18282] + MEM[18690];
assign MEM[27604] = MEM[18283] + MEM[19044];
assign MEM[27605] = MEM[18285] + MEM[18469];
assign MEM[27606] = MEM[18288] + MEM[18865];
assign MEM[27607] = MEM[18289] + MEM[18648];
assign MEM[27608] = MEM[18290] + MEM[18807];
assign MEM[27609] = MEM[18292] + MEM[19241];
assign MEM[27610] = MEM[18293] + MEM[18836];
assign MEM[27611] = MEM[18295] + MEM[18511];
assign MEM[27612] = MEM[18296] + MEM[18475];
assign MEM[27613] = MEM[18297] + MEM[18514];
assign MEM[27614] = MEM[18306] + MEM[18354];
assign MEM[27615] = MEM[18310] + MEM[18395];
assign MEM[27616] = MEM[18313] + MEM[18496];
assign MEM[27617] = MEM[18317] + MEM[18701];
assign MEM[27618] = MEM[18324] + MEM[18918];
assign MEM[27619] = MEM[18326] + MEM[18346];
assign MEM[27620] = MEM[18327] + MEM[18528];
assign MEM[27621] = MEM[18328] + MEM[18509];
assign MEM[27622] = MEM[18330] + MEM[18809];
assign MEM[27623] = MEM[18331] + MEM[18411];
assign MEM[27624] = MEM[18335] + MEM[18644];
assign MEM[27625] = MEM[18337] + MEM[18837];
assign MEM[27626] = MEM[18339] + MEM[18618];
assign MEM[27627] = MEM[18341] + MEM[19068];
assign MEM[27628] = MEM[18348] + MEM[18540];
assign MEM[27629] = MEM[18349] + MEM[19100];
assign MEM[27630] = MEM[18351] + MEM[18937];
assign MEM[27631] = MEM[18365] + MEM[19458];
assign MEM[27632] = MEM[18366] + MEM[18383];
assign MEM[27633] = MEM[18368] + MEM[19186];
assign MEM[27634] = MEM[18371] + MEM[18546];
assign MEM[27635] = MEM[18376] + MEM[19306];
assign MEM[27636] = MEM[18377] + MEM[18944];
assign MEM[27637] = MEM[18380] + MEM[18449];
assign MEM[27638] = MEM[18386] + MEM[19185];
assign MEM[27639] = MEM[18392] + MEM[18737];
assign MEM[27640] = MEM[18393] + MEM[18425];
assign MEM[27641] = MEM[18394] + MEM[18658];
assign MEM[27642] = MEM[18396] + MEM[18544];
assign MEM[27643] = MEM[18399] + MEM[18525];
assign MEM[27644] = MEM[18403] + MEM[18450];
assign MEM[27645] = MEM[18409] + MEM[18497];
assign MEM[27646] = MEM[18410] + MEM[18468];
assign MEM[27647] = MEM[18412] + MEM[18506];
assign MEM[27648] = MEM[18414] + MEM[18829];
assign MEM[27649] = MEM[18415] + MEM[19175];
assign MEM[27650] = MEM[18416] + MEM[18650];
assign MEM[27651] = MEM[18417] + MEM[18577];
assign MEM[27652] = MEM[18418] + MEM[18850];
assign MEM[27653] = MEM[18419] + MEM[18428];
assign MEM[27654] = MEM[18420] + MEM[18588];
assign MEM[27655] = MEM[18421] + MEM[19041];
assign MEM[27656] = MEM[18422] + MEM[18982];
assign MEM[27657] = MEM[18423] + MEM[18845];
assign MEM[27658] = MEM[18427] + MEM[18685];
assign MEM[27659] = MEM[18430] + MEM[19383];
assign MEM[27660] = MEM[18432] + MEM[18578];
assign MEM[27661] = MEM[18439] + MEM[18782];
assign MEM[27662] = MEM[18443] + MEM[18909];
assign MEM[27663] = MEM[18448] + MEM[19348];
assign MEM[27664] = MEM[18455] + MEM[18858];
assign MEM[27665] = MEM[18459] + MEM[18980];
assign MEM[27666] = MEM[18460] + MEM[18548];
assign MEM[27667] = MEM[18465] + MEM[18914];
assign MEM[27668] = MEM[18466] + MEM[18900];
assign MEM[27669] = MEM[18470] + MEM[18869];
assign MEM[27670] = MEM[18471] + MEM[19173];
assign MEM[27671] = MEM[18479] + MEM[18513];
assign MEM[27672] = MEM[18486] + MEM[19315];
assign MEM[27673] = MEM[18488] + MEM[18818];
assign MEM[27674] = MEM[18489] + MEM[18704];
assign MEM[27675] = MEM[18493] + MEM[19723];
assign MEM[27676] = MEM[18499] + MEM[18670];
assign MEM[27677] = MEM[18504] + MEM[18695];
assign MEM[27678] = MEM[18508] + MEM[19467];
assign MEM[27679] = MEM[18512] + MEM[18633];
assign MEM[27680] = MEM[18519] + MEM[18743];
assign MEM[27681] = MEM[18524] + MEM[19001];
assign MEM[27682] = MEM[18527] + MEM[18791];
assign MEM[27683] = MEM[18529] + MEM[18744];
assign MEM[27684] = MEM[18530] + MEM[18612];
assign MEM[27685] = MEM[18531] + MEM[19113];
assign MEM[27686] = MEM[18534] + MEM[18904];
assign MEM[27687] = MEM[18538] + MEM[19013];
assign MEM[27688] = MEM[18541] + MEM[18749];
assign MEM[27689] = MEM[18542] + MEM[18770];
assign MEM[27690] = MEM[18543] + MEM[18678];
assign MEM[27691] = MEM[18547] + MEM[18781];
assign MEM[27692] = MEM[18550] + MEM[19197];
assign MEM[27693] = MEM[18551] + MEM[19373];
assign MEM[27694] = MEM[18553] + MEM[18560];
assign MEM[27695] = MEM[18562] + MEM[19097];
assign MEM[27696] = MEM[18565] + MEM[19057];
assign MEM[27697] = MEM[18571] + MEM[18719];
assign MEM[27698] = MEM[18572] + MEM[18703];
assign MEM[27699] = MEM[18574] + MEM[18765];
assign MEM[27700] = MEM[18582] + MEM[18957];
assign MEM[27701] = MEM[18584] + MEM[18754];
assign MEM[27702] = MEM[18585] + MEM[19129];
assign MEM[27703] = MEM[18586] + MEM[18823];
assign MEM[27704] = MEM[18589] + MEM[19499];
assign MEM[27705] = MEM[18594] + MEM[18645];
assign MEM[27706] = MEM[18595] + MEM[19014];
assign MEM[27707] = MEM[18597] + MEM[19286];
assign MEM[27708] = MEM[18600] + MEM[18713];
assign MEM[27709] = MEM[18605] + MEM[18683];
assign MEM[27710] = MEM[18611] + MEM[19258];
assign MEM[27711] = MEM[18614] + MEM[18705];
assign MEM[27712] = MEM[18624] + MEM[19027];
assign MEM[27713] = MEM[18626] + MEM[18752];
assign MEM[27714] = MEM[18627] + MEM[18654];
assign MEM[27715] = MEM[18628] + MEM[18901];
assign MEM[27716] = MEM[18630] + MEM[18978];
assign MEM[27717] = MEM[18631] + MEM[18859];
assign MEM[27718] = MEM[18632] + MEM[18709];
assign MEM[27719] = MEM[18634] + MEM[18647];
assign MEM[27720] = MEM[18637] + MEM[18889];
assign MEM[27721] = MEM[18638] + MEM[18821];
assign MEM[27722] = MEM[18639] + MEM[18831];
assign MEM[27723] = MEM[18641] + MEM[19220];
assign MEM[27724] = MEM[18642] + MEM[18787];
assign MEM[27725] = MEM[18649] + MEM[18848];
assign MEM[27726] = MEM[18651] + MEM[18851];
assign MEM[27727] = MEM[18653] + MEM[19732];
assign MEM[27728] = MEM[18656] + MEM[19018];
assign MEM[27729] = MEM[18659] + MEM[18665];
assign MEM[27730] = MEM[18661] + MEM[19004];
assign MEM[27731] = MEM[18666] + MEM[19240];
assign MEM[27732] = MEM[18668] + MEM[18890];
assign MEM[27733] = MEM[18671] + MEM[18996];
assign MEM[27734] = MEM[18673] + MEM[18860];
assign MEM[27735] = MEM[18675] + MEM[19243];
assign MEM[27736] = MEM[18676] + MEM[18857];
assign MEM[27737] = MEM[18677] + MEM[18943];
assign MEM[27738] = MEM[18681] + MEM[19167];
assign MEM[27739] = MEM[18686] + MEM[19043];
assign MEM[27740] = MEM[18692] + MEM[19257];
assign MEM[27741] = MEM[18697] + MEM[19881];
assign MEM[27742] = MEM[18698] + MEM[19077];
assign MEM[27743] = MEM[18699] + MEM[18949];
assign MEM[27744] = MEM[18707] + MEM[19300];
assign MEM[27745] = MEM[18710] + MEM[18835];
assign MEM[27746] = MEM[18711] + MEM[18897];
assign MEM[27747] = MEM[18714] + MEM[19385];
assign MEM[27748] = MEM[18720] + MEM[19529];
assign MEM[27749] = MEM[18723] + MEM[18853];
assign MEM[27750] = MEM[18724] + MEM[19546];
assign MEM[27751] = MEM[18725] + MEM[18838];
assign MEM[27752] = MEM[18727] + MEM[19267];
assign MEM[27753] = MEM[18728] + MEM[19063];
assign MEM[27754] = MEM[18731] + MEM[18894];
assign MEM[27755] = MEM[18734] + MEM[18867];
assign MEM[27756] = MEM[18739] + MEM[18847];
assign MEM[27757] = MEM[18746] + MEM[19951];
assign MEM[27758] = MEM[18747] + MEM[18878];
assign MEM[27759] = MEM[18748] + MEM[19122];
assign MEM[27760] = MEM[18750] + MEM[18929];
assign MEM[27761] = MEM[18751] + MEM[18990];
assign MEM[27762] = MEM[18753] + MEM[19158];
assign MEM[27763] = MEM[18756] + MEM[19309];
assign MEM[27764] = MEM[18759] + MEM[18806];
assign MEM[27765] = MEM[18760] + MEM[19493];
assign MEM[27766] = MEM[18761] + MEM[19109];
assign MEM[27767] = MEM[18764] + MEM[18768];
assign MEM[27768] = MEM[18767] + MEM[19007];
assign MEM[27769] = MEM[18769] + MEM[18783];
assign MEM[27770] = MEM[18775] + MEM[18969];
assign MEM[27771] = MEM[18776] + MEM[18947];
assign MEM[27772] = MEM[18778] + MEM[20273];
assign MEM[27773] = MEM[18779] + MEM[18801];
assign MEM[27774] = MEM[18788] + MEM[19107];
assign MEM[27775] = MEM[18792] + MEM[19314];
assign MEM[27776] = MEM[18794] + MEM[18922];
assign MEM[27777] = MEM[18797] + MEM[19123];
assign MEM[27778] = MEM[18798] + MEM[18910];
assign MEM[27779] = MEM[18803] + MEM[19363];
assign MEM[27780] = MEM[18805] + MEM[19151];
assign MEM[27781] = MEM[18808] + MEM[18874];
assign MEM[27782] = MEM[18812] + MEM[19132];
assign MEM[27783] = MEM[18814] + MEM[18953];
assign MEM[27784] = MEM[18820] + MEM[19390];
assign MEM[27785] = MEM[18822] + MEM[19460];
assign MEM[27786] = MEM[18826] + MEM[19066];
assign MEM[27787] = MEM[18827] + MEM[19364];
assign MEM[27788] = MEM[18828] + MEM[19020];
assign MEM[27789] = MEM[18830] + MEM[19073];
assign MEM[27790] = MEM[18832] + MEM[19433];
assign MEM[27791] = MEM[18834] + MEM[19844];
assign MEM[27792] = MEM[18843] + MEM[18971];
assign MEM[27793] = MEM[18844] + MEM[20047];
assign MEM[27794] = MEM[18861] + MEM[19607];
assign MEM[27795] = MEM[18862] + MEM[19251];
assign MEM[27796] = MEM[18864] + MEM[18989];
assign MEM[27797] = MEM[18866] + MEM[19766];
assign MEM[27798] = MEM[18870] + MEM[19224];
assign MEM[27799] = MEM[18873] + MEM[19191];
assign MEM[27800] = MEM[18876] + MEM[18951];
assign MEM[27801] = MEM[18877] + MEM[19430];
assign MEM[27802] = MEM[18880] + MEM[19252];
assign MEM[27803] = MEM[18881] + MEM[19278];
assign MEM[27804] = MEM[18882] + MEM[19368];
assign MEM[27805] = MEM[18883] + MEM[18892];
assign MEM[27806] = MEM[18884] + MEM[19418];
assign MEM[27807] = MEM[18893] + MEM[19636];
assign MEM[27808] = MEM[18898] + MEM[19571];
assign MEM[27809] = MEM[18906] + MEM[19035];
assign MEM[27810] = MEM[18907] + MEM[19938];
assign MEM[27811] = MEM[18908] + MEM[19423];
assign MEM[27812] = MEM[18912] + MEM[19866];
assign MEM[27813] = MEM[18920] + MEM[19369];
assign MEM[27814] = MEM[18923] + MEM[19023];
assign MEM[27815] = MEM[18924] + MEM[19103];
assign MEM[27816] = MEM[18925] + MEM[20063];
assign MEM[27817] = MEM[18928] + MEM[19464];
assign MEM[27818] = MEM[18932] + MEM[18968];
assign MEM[27819] = MEM[18933] + MEM[19536];
assign MEM[27820] = MEM[18934] + MEM[19207];
assign MEM[27821] = MEM[18938] + MEM[19254];
assign MEM[27822] = MEM[18939] + MEM[19169];
assign MEM[27823] = MEM[18940] + MEM[19166];
assign MEM[27824] = MEM[18950] + MEM[19052];
assign MEM[27825] = MEM[18952] + MEM[19235];
assign MEM[27826] = MEM[18954] + MEM[19993];
assign MEM[27827] = MEM[18955] + MEM[19223];
assign MEM[27828] = MEM[18959] + MEM[18960];
assign MEM[27829] = MEM[18963] + MEM[19233];
assign MEM[27830] = MEM[18964] + MEM[19048];
assign MEM[27831] = MEM[18965] + MEM[19814];
assign MEM[27832] = MEM[18973] + MEM[19810];
assign MEM[27833] = MEM[18974] + MEM[19088];
assign MEM[27834] = MEM[18981] + MEM[19124];
assign MEM[27835] = MEM[18983] + MEM[19279];
assign MEM[27836] = MEM[18984] + MEM[19709];
assign MEM[27837] = MEM[18986] + MEM[19795];
assign MEM[27838] = MEM[18988] + MEM[19105];
assign MEM[27839] = MEM[18993] + MEM[19070];
assign MEM[27840] = MEM[18994] + MEM[19011];
assign MEM[27841] = MEM[18997] + MEM[19053];
assign MEM[27842] = MEM[19000] + MEM[19519];
assign MEM[27843] = MEM[19002] + MEM[19111];
assign MEM[27844] = MEM[19003] + MEM[19212];
assign MEM[27845] = MEM[19006] + MEM[19112];
assign MEM[27846] = MEM[19012] + MEM[19160];
assign MEM[27847] = MEM[19016] + MEM[19294];
assign MEM[27848] = MEM[19022] + MEM[19104];
assign MEM[27849] = MEM[19024] + MEM[19513];
assign MEM[27850] = MEM[19025] + MEM[19290];
assign MEM[27851] = MEM[19026] + MEM[19457];
assign MEM[27852] = MEM[19028] + MEM[19106];
assign MEM[27853] = MEM[19031] + MEM[19461];
assign MEM[27854] = MEM[19032] + MEM[19377];
assign MEM[27855] = MEM[19033] + MEM[19505];
assign MEM[27856] = MEM[19036] + MEM[19358];
assign MEM[27857] = MEM[19037] + MEM[19065];
assign MEM[27858] = MEM[19038] + MEM[19163];
assign MEM[27859] = MEM[19039] + MEM[19990];
assign MEM[27860] = MEM[19042] + MEM[19451];
assign MEM[27861] = MEM[19046] + MEM[19284];
assign MEM[27862] = MEM[19047] + MEM[19454];
assign MEM[27863] = MEM[19049] + MEM[19146];
assign MEM[27864] = MEM[19050] + MEM[19353];
assign MEM[27865] = MEM[19055] + MEM[19572];
assign MEM[27866] = MEM[19056] + MEM[19532];
assign MEM[27867] = MEM[19058] + MEM[19453];
assign MEM[27868] = MEM[19060] + MEM[19208];
assign MEM[27869] = MEM[19062] + MEM[19142];
assign MEM[27870] = MEM[19064] + MEM[19537];
assign MEM[27871] = MEM[19067] + MEM[20255];
assign MEM[27872] = MEM[19069] + MEM[20114];
assign MEM[27873] = MEM[19071] + MEM[20846];
assign MEM[27874] = MEM[19074] + MEM[19644];
assign MEM[27875] = MEM[19078] + MEM[19804];
assign MEM[27876] = MEM[19079] + MEM[19318];
assign MEM[27877] = MEM[19084] + MEM[19301];
assign MEM[27878] = MEM[19086] + MEM[19248];
assign MEM[27879] = MEM[19087] + MEM[19255];
assign MEM[27880] = MEM[19090] + MEM[19658];
assign MEM[27881] = MEM[19092] + MEM[19590];
assign MEM[27882] = MEM[19093] + MEM[19346];
assign MEM[27883] = MEM[19094] + MEM[19230];
assign MEM[27884] = MEM[19095] + MEM[19728];
assign MEM[27885] = MEM[19102] + MEM[19205];
assign MEM[27886] = MEM[19110] + MEM[19631];
assign MEM[27887] = MEM[19117] + MEM[19873];
assign MEM[27888] = MEM[19118] + MEM[20129];
assign MEM[27889] = MEM[19119] + MEM[19594];
assign MEM[27890] = MEM[19120] + MEM[19136];
assign MEM[27891] = MEM[19126] + MEM[19326];
assign MEM[27892] = MEM[19128] + MEM[19388];
assign MEM[27893] = MEM[19131] + MEM[19362];
assign MEM[27894] = MEM[19133] + MEM[19189];
assign MEM[27895] = MEM[19135] + MEM[19216];
assign MEM[27896] = MEM[19139] + MEM[20040];
assign MEM[27897] = MEM[19141] + MEM[19442];
assign MEM[27898] = MEM[19145] + MEM[19264];
assign MEM[27899] = MEM[19147] + MEM[19500];
assign MEM[27900] = MEM[19148] + MEM[19149];
assign MEM[27901] = MEM[19153] + MEM[19913];
assign MEM[27902] = MEM[19154] + MEM[19161];
assign MEM[27903] = MEM[19156] + MEM[19209];
assign MEM[27904] = MEM[19157] + MEM[19198];
assign MEM[27905] = MEM[19162] + MEM[19633];
assign MEM[27906] = MEM[19168] + MEM[19730];
assign MEM[27907] = MEM[19170] + MEM[19496];
assign MEM[27908] = MEM[19172] + MEM[19717];
assign MEM[27909] = MEM[19174] + MEM[19488];
assign MEM[27910] = MEM[19179] + MEM[19180];
assign MEM[27911] = MEM[19181] + MEM[19969];
assign MEM[27912] = MEM[19182] + MEM[19557];
assign MEM[27913] = MEM[19184] + MEM[19725];
assign MEM[27914] = MEM[19187] + MEM[19389];
assign MEM[27915] = MEM[19190] + MEM[19345];
assign MEM[27916] = MEM[19192] + MEM[19510];
assign MEM[27917] = MEM[19193] + MEM[19824];
assign MEM[27918] = MEM[19195] + MEM[19931];
assign MEM[27919] = MEM[19196] + MEM[19923];
assign MEM[27920] = MEM[19202] + MEM[19269];
assign MEM[27921] = MEM[19204] + MEM[19731];
assign MEM[27922] = MEM[19206] + MEM[19776];
assign MEM[27923] = MEM[19210] + MEM[19404];
assign MEM[27924] = MEM[19213] + MEM[19411];
assign MEM[27925] = MEM[19215] + MEM[19288];
assign MEM[27926] = MEM[19217] + MEM[19394];
assign MEM[27927] = MEM[19218] + MEM[19476];
assign MEM[27928] = MEM[19219] + MEM[19285];
assign MEM[27929] = MEM[19221] + MEM[19697];
assign MEM[27930] = MEM[19222] + MEM[19919];
assign MEM[27931] = MEM[19229] + MEM[19324];
assign MEM[27932] = MEM[19231] + MEM[20937];
assign MEM[27933] = MEM[19232] + MEM[19474];
assign MEM[27934] = MEM[19234] + MEM[19397];
assign MEM[27935] = MEM[19237] + MEM[20160];
assign MEM[27936] = MEM[19238] + MEM[19400];
assign MEM[27937] = MEM[19245] + MEM[19986];
assign MEM[27938] = MEM[19246] + MEM[19507];
assign MEM[27939] = MEM[19249] + MEM[19889];
assign MEM[27940] = MEM[19253] + MEM[19405];
assign MEM[27941] = MEM[19256] + MEM[20368];
assign MEM[27942] = MEM[19259] + MEM[19365];
assign MEM[27943] = MEM[19261] + MEM[19281];
assign MEM[27944] = MEM[19262] + MEM[19349];
assign MEM[27945] = MEM[19265] + MEM[19490];
assign MEM[27946] = MEM[19268] + MEM[20011];
assign MEM[27947] = MEM[19270] + MEM[19305];
assign MEM[27948] = MEM[19272] + MEM[20180];
assign MEM[27949] = MEM[19273] + MEM[19356];
assign MEM[27950] = MEM[19274] + MEM[19440];
assign MEM[27951] = MEM[19277] + MEM[19784];
assign MEM[27952] = MEM[19280] + MEM[19292];
assign MEM[27953] = MEM[19287] + MEM[19379];
assign MEM[27954] = MEM[19289] + MEM[19325];
assign MEM[27955] = MEM[19291] + MEM[19443];
assign MEM[27956] = MEM[19293] + MEM[19503];
assign MEM[27957] = MEM[19298] + MEM[19331];
assign MEM[27958] = MEM[19299] + MEM[19611];
assign MEM[27959] = MEM[19302] + MEM[19313];
assign MEM[27960] = MEM[19303] + MEM[19387];
assign MEM[27961] = MEM[19307] + MEM[19334];
assign MEM[27962] = MEM[19310] + MEM[19605];
assign MEM[27963] = MEM[19311] + MEM[19321];
assign MEM[27964] = MEM[19312] + MEM[19929];
assign MEM[27965] = MEM[19316] + MEM[20198];
assign MEM[27966] = MEM[19322] + MEM[19542];
assign MEM[27967] = MEM[19323] + MEM[19699];
assign MEM[27968] = MEM[19327] + MEM[19854];
assign MEM[27969] = MEM[19328] + MEM[19909];
assign MEM[27970] = MEM[19329] + MEM[19465];
assign MEM[27971] = MEM[19330] + MEM[19455];
assign MEM[27972] = MEM[19332] + MEM[19447];
assign MEM[27973] = MEM[19333] + MEM[19643];
assign MEM[27974] = MEM[19335] + MEM[19541];
assign MEM[27975] = MEM[19337] + MEM[19339];
assign MEM[27976] = MEM[19338] + MEM[19562];
assign MEM[27977] = MEM[19340] + MEM[19692];
assign MEM[27978] = MEM[19344] + MEM[19991];
assign MEM[27979] = MEM[19347] + MEM[19822];
assign MEM[27980] = MEM[19350] + MEM[19498];
assign MEM[27981] = MEM[19351] + MEM[19452];
assign MEM[27982] = MEM[19352] + MEM[19680];
assign MEM[27983] = MEM[19354] + MEM[19361];
assign MEM[27984] = MEM[19360] + MEM[19580];
assign MEM[27985] = MEM[19366] + MEM[19729];
assign MEM[27986] = MEM[19367] + MEM[19626];
assign MEM[27987] = MEM[19370] + MEM[19592];
assign MEM[27988] = MEM[19372] + MEM[19879];
assign MEM[27989] = MEM[19374] + MEM[19805];
assign MEM[27990] = MEM[19375] + MEM[20301];
assign MEM[27991] = MEM[19378] + MEM[19762];
assign MEM[27992] = MEM[19380] + MEM[19509];
assign MEM[27993] = MEM[19386] + MEM[20661];
assign MEM[27994] = MEM[19391] + MEM[19597];
assign MEM[27995] = MEM[19392] + MEM[20623];
assign MEM[27996] = MEM[19396] + MEM[19883];
assign MEM[27997] = MEM[19398] + MEM[19494];
assign MEM[27998] = MEM[19401] + MEM[19504];
assign MEM[27999] = MEM[19402] + MEM[19586];
assign MEM[28000] = MEM[19406] + MEM[19610];
assign MEM[28001] = MEM[19407] + MEM[20427];
assign MEM[28002] = MEM[19408] + MEM[19525];
assign MEM[28003] = MEM[19410] + MEM[19685];
assign MEM[28004] = MEM[19413] + MEM[19973];
assign MEM[28005] = MEM[19417] + MEM[20092];
assign MEM[28006] = MEM[19420] + MEM[19778];
assign MEM[28007] = MEM[19421] + MEM[19899];
assign MEM[28008] = MEM[19422] + MEM[19591];
assign MEM[28009] = MEM[19424] + MEM[19574];
assign MEM[28010] = MEM[19426] + MEM[19813];
assign MEM[28011] = MEM[19427] + MEM[20045];
assign MEM[28012] = MEM[19428] + MEM[21369];
assign MEM[28013] = MEM[19429] + MEM[19563];
assign MEM[28014] = MEM[19432] + MEM[20000];
assign MEM[28015] = MEM[19435] + MEM[19927];
assign MEM[28016] = MEM[19436] + MEM[19466];
assign MEM[28017] = MEM[19438] + MEM[20291];
assign MEM[28018] = MEM[19444] + MEM[19472];
assign MEM[28019] = MEM[19446] + MEM[19514];
assign MEM[28020] = MEM[19448] + MEM[20420];
assign MEM[28021] = MEM[19449] + MEM[19534];
assign MEM[28022] = MEM[19450] + MEM[19742];
assign MEM[28023] = MEM[19456] + MEM[19601];
assign MEM[28024] = MEM[19459] + MEM[19629];
assign MEM[28025] = MEM[19462] + MEM[19696];
assign MEM[28026] = MEM[19468] + MEM[19704];
assign MEM[28027] = MEM[19469] + MEM[19695];
assign MEM[28028] = MEM[19470] + MEM[20014];
assign MEM[28029] = MEM[19471] + MEM[19847];
assign MEM[28030] = MEM[19473] + MEM[19819];
assign MEM[28031] = MEM[19475] + MEM[19833];
assign MEM[28032] = MEM[19477] + MEM[19647];
assign MEM[28033] = MEM[19480] + MEM[19829];
assign MEM[28034] = MEM[19484] + MEM[20001];
assign MEM[28035] = MEM[19486] + MEM[20106];
assign MEM[28036] = MEM[19489] + MEM[19734];
assign MEM[28037] = MEM[19492] + MEM[19664];
assign MEM[28038] = MEM[19495] + MEM[19746];
assign MEM[28039] = MEM[19502] + MEM[20064];
assign MEM[28040] = MEM[19506] + MEM[19985];
assign MEM[28041] = MEM[19508] + MEM[19958];
assign MEM[28042] = MEM[19511] + MEM[19589];
assign MEM[28043] = MEM[19515] + MEM[19568];
assign MEM[28044] = MEM[19516] + MEM[19890];
assign MEM[28045] = MEM[19517] + MEM[19957];
assign MEM[28046] = MEM[19518] + MEM[19910];
assign MEM[28047] = MEM[19520] + MEM[19635];
assign MEM[28048] = MEM[19522] + MEM[19553];
assign MEM[28049] = MEM[19523] + MEM[19808];
assign MEM[28050] = MEM[19524] + MEM[19920];
assign MEM[28051] = MEM[19526] + MEM[20055];
assign MEM[28052] = MEM[19527] + MEM[19552];
assign MEM[28053] = MEM[19528] + MEM[20300];
assign MEM[28054] = MEM[19530] + MEM[19727];
assign MEM[28055] = MEM[19531] + MEM[19670];
assign MEM[28056] = MEM[19533] + MEM[19780];
assign MEM[28057] = MEM[19538] + MEM[19615];
assign MEM[28058] = MEM[19539] + MEM[20051];
assign MEM[28059] = MEM[19540] + MEM[20013];
assign MEM[28060] = MEM[19543] + MEM[20006];
assign MEM[28061] = MEM[19544] + MEM[20208];
assign MEM[28062] = MEM[19547] + MEM[19548];
assign MEM[28063] = MEM[19549] + MEM[20386];
assign MEM[28064] = MEM[19550] + MEM[20034];
assign MEM[28065] = MEM[19551] + MEM[20058];
assign MEM[28066] = MEM[19555] + MEM[19785];
assign MEM[28067] = MEM[19559] + MEM[19686];
assign MEM[28068] = MEM[19560] + MEM[19718];
assign MEM[28069] = MEM[19561] + MEM[20117];
assign MEM[28070] = MEM[19567] + MEM[19584];
assign MEM[28071] = MEM[19569] + MEM[20178];
assign MEM[28072] = MEM[19570] + MEM[20070];
assign MEM[28073] = MEM[19576] + MEM[19756];
assign MEM[28074] = MEM[19577] + MEM[19836];
assign MEM[28075] = MEM[19578] + MEM[20514];
assign MEM[28076] = MEM[19581] + MEM[19671];
assign MEM[28077] = MEM[19582] + MEM[19740];
assign MEM[28078] = MEM[19583] + MEM[19621];
assign MEM[28079] = MEM[19587] + MEM[19858];
assign MEM[28080] = MEM[19593] + MEM[20107];
assign MEM[28081] = MEM[19595] + MEM[20078];
assign MEM[28082] = MEM[19598] + MEM[20350];
assign MEM[28083] = MEM[19599] + MEM[20138];
assign MEM[28084] = MEM[19602] + MEM[19733];
assign MEM[28085] = MEM[19603] + MEM[19632];
assign MEM[28086] = MEM[19606] + MEM[19863];
assign MEM[28087] = MEM[19609] + MEM[19668];
assign MEM[28088] = MEM[19612] + MEM[19980];
assign MEM[28089] = MEM[19613] + MEM[19678];
assign MEM[28090] = MEM[19614] + MEM[19790];
assign MEM[28091] = MEM[19616] + MEM[19763];
assign MEM[28092] = MEM[19619] + MEM[19679];
assign MEM[28093] = MEM[19620] + MEM[19758];
assign MEM[28094] = MEM[19622] + MEM[19684];
assign MEM[28095] = MEM[19624] + MEM[20050];
assign MEM[28096] = MEM[19625] + MEM[19650];
assign MEM[28097] = MEM[19627] + MEM[19774];
assign MEM[28098] = MEM[19630] + MEM[19867];
assign MEM[28099] = MEM[19634] + MEM[20203];
assign MEM[28100] = MEM[19640] + MEM[19924];
assign MEM[28101] = MEM[19641] + MEM[19651];
assign MEM[28102] = MEM[19646] + MEM[19936];
assign MEM[28103] = MEM[19648] + MEM[20049];
assign MEM[28104] = MEM[19649] + MEM[19974];
assign MEM[28105] = MEM[19652] + MEM[20200];
assign MEM[28106] = MEM[19653] + MEM[19964];
assign MEM[28107] = MEM[19654] + MEM[19870];
assign MEM[28108] = MEM[19655] + MEM[20286];
assign MEM[28109] = MEM[19657] + MEM[20086];
assign MEM[28110] = MEM[19660] + MEM[19802];
assign MEM[28111] = MEM[19661] + MEM[19967];
assign MEM[28112] = MEM[19662] + MEM[19767];
assign MEM[28113] = MEM[19663] + MEM[19976];
assign MEM[28114] = MEM[19665] + MEM[20399];
assign MEM[28115] = MEM[19666] + MEM[20018];
assign MEM[28116] = MEM[19673] + MEM[19988];
assign MEM[28117] = MEM[19674] + MEM[20632];
assign MEM[28118] = MEM[19675] + MEM[20384];
assign MEM[28119] = MEM[19676] + MEM[20223];
assign MEM[28120] = MEM[19681] + MEM[19892];
assign MEM[28121] = MEM[19682] + MEM[20400];
assign MEM[28122] = MEM[19683] + MEM[20023];
assign MEM[28123] = MEM[19687] + MEM[19741];
assign MEM[28124] = MEM[19688] + MEM[19897];
assign MEM[28125] = MEM[19698] + MEM[19989];
assign MEM[28126] = MEM[19701] + MEM[20769];
assign MEM[28127] = MEM[19702] + MEM[19736];
assign MEM[28128] = MEM[19703] + MEM[20490];
assign MEM[28129] = MEM[19707] + MEM[19995];
assign MEM[28130] = MEM[19708] + MEM[19753];
assign MEM[28131] = MEM[19712] + MEM[20569];
assign MEM[28132] = MEM[19714] + MEM[19772];
assign MEM[28133] = MEM[19715] + MEM[19748];
assign MEM[28134] = MEM[19716] + MEM[20141];
assign MEM[28135] = MEM[19719] + MEM[19877];
assign MEM[28136] = MEM[19726] + MEM[20083];
assign MEM[28137] = MEM[19735] + MEM[19862];
assign MEM[28138] = MEM[19737] + MEM[20191];
assign MEM[28139] = MEM[19738] + MEM[19747];
assign MEM[28140] = MEM[19744] + MEM[20270];
assign MEM[28141] = MEM[19745] + MEM[19885];
assign MEM[28142] = MEM[19749] + MEM[20169];
assign MEM[28143] = MEM[19750] + MEM[20062];
assign MEM[28144] = MEM[19751] + MEM[20523];
assign MEM[28145] = MEM[19752] + MEM[20394];
assign MEM[28146] = MEM[19757] + MEM[20532];
assign MEM[28147] = MEM[19760] + MEM[20137];
assign MEM[28148] = MEM[19761] + MEM[20268];
assign MEM[28149] = MEM[19768] + MEM[19955];
assign MEM[28150] = MEM[19769] + MEM[20101];
assign MEM[28151] = MEM[19770] + MEM[20094];
assign MEM[28152] = MEM[19773] + MEM[20447];
assign MEM[28153] = MEM[19775] + MEM[19917];
assign MEM[28154] = MEM[19779] + MEM[19834];
assign MEM[28155] = MEM[19781] + MEM[20104];
assign MEM[28156] = MEM[19782] + MEM[19872];
assign MEM[28157] = MEM[19783] + MEM[20087];
assign MEM[28158] = MEM[19786] + MEM[20486];
assign MEM[28159] = MEM[19791] + MEM[19842];
assign MEM[28160] = MEM[19792] + MEM[20329];
assign MEM[28161] = MEM[19793] + MEM[19830];
assign MEM[28162] = MEM[19794] + MEM[19904];
assign MEM[28163] = MEM[19797] + MEM[19887];
assign MEM[28164] = MEM[19798] + MEM[19871];
assign MEM[28165] = MEM[19809] + MEM[19839];
assign MEM[28166] = MEM[19812] + MEM[19826];
assign MEM[28167] = MEM[19815] + MEM[19898];
assign MEM[28168] = MEM[19816] + MEM[19978];
assign MEM[28169] = MEM[19817] + MEM[19960];
assign MEM[28170] = MEM[19818] + MEM[20163];
assign MEM[28171] = MEM[19820] + MEM[20100];
assign MEM[28172] = MEM[19825] + MEM[19903];
assign MEM[28173] = MEM[19831] + MEM[20287];
assign MEM[28174] = MEM[19840] + MEM[19922];
assign MEM[28175] = MEM[19841] + MEM[19930];
assign MEM[28176] = MEM[19845] + MEM[20004];
assign MEM[28177] = MEM[19849] + MEM[19875];
assign MEM[28178] = MEM[19850] + MEM[20182];
assign MEM[28179] = MEM[19851] + MEM[20032];
assign MEM[28180] = MEM[19852] + MEM[20119];
assign MEM[28181] = MEM[19853] + MEM[20152];
assign MEM[28182] = MEM[19855] + MEM[20283];
assign MEM[28183] = MEM[19857] + MEM[20019];
assign MEM[28184] = MEM[19859] + MEM[20103];
assign MEM[28185] = MEM[19860] + MEM[20635];
assign MEM[28186] = MEM[19861] + MEM[20190];
assign MEM[28187] = MEM[19864] + MEM[20136];
assign MEM[28188] = MEM[19868] + MEM[20312];
assign MEM[28189] = MEM[19869] + MEM[20426];
assign MEM[28190] = MEM[19874] + MEM[19888];
assign MEM[28191] = MEM[19876] + MEM[21121];
assign MEM[28192] = MEM[19882] + MEM[20611];
assign MEM[28193] = MEM[19884] + MEM[20036];
assign MEM[28194] = MEM[19893] + MEM[20009];
assign MEM[28195] = MEM[19894] + MEM[20108];
assign MEM[28196] = MEM[19896] + MEM[20041];
assign MEM[28197] = MEM[19901] + MEM[19912];
assign MEM[28198] = MEM[19905] + MEM[20253];
assign MEM[28199] = MEM[19906] + MEM[19968];
assign MEM[28200] = MEM[19907] + MEM[19983];
assign MEM[28201] = MEM[19908] + MEM[20409];
assign MEM[28202] = MEM[19914] + MEM[20474];
assign MEM[28203] = MEM[19918] + MEM[20081];
assign MEM[28204] = MEM[19921] + MEM[20258];
assign MEM[28205] = MEM[19925] + MEM[20197];
assign MEM[28206] = MEM[19928] + MEM[20266];
assign MEM[28207] = MEM[19932] + MEM[19952];
assign MEM[28208] = MEM[19933] + MEM[19965];
assign MEM[28209] = MEM[19934] + MEM[20463];
assign MEM[28210] = MEM[19935] + MEM[20282];
assign MEM[28211] = MEM[19937] + MEM[20020];
assign MEM[28212] = MEM[19939] + MEM[20348];
assign MEM[28213] = MEM[19940] + MEM[20476];
assign MEM[28214] = MEM[19941] + MEM[20044];
assign MEM[28215] = MEM[19942] + MEM[20904];
assign MEM[28216] = MEM[19943] + MEM[20121];
assign MEM[28217] = MEM[19944] + MEM[20128];
assign MEM[28218] = MEM[19945] + MEM[19970];
assign MEM[28219] = MEM[19946] + MEM[20142];
assign MEM[28220] = MEM[19947] + MEM[20167];
assign MEM[28221] = MEM[19949] + MEM[20374];
assign MEM[28222] = MEM[19953] + MEM[20252];
assign MEM[28223] = MEM[19954] + MEM[20015];
assign MEM[28224] = MEM[19959] + MEM[20589];
assign MEM[28225] = MEM[19962] + MEM[20185];
assign MEM[28226] = MEM[19963] + MEM[20930];
assign MEM[28227] = MEM[19966] + MEM[20387];
assign MEM[28228] = MEM[19971] + MEM[20111];
assign MEM[28229] = MEM[19975] + MEM[20284];
assign MEM[28230] = MEM[19977] + MEM[20037];
assign MEM[28231] = MEM[19979] + MEM[20362];
assign MEM[28232] = MEM[19981] + MEM[20161];
assign MEM[28233] = MEM[19982] + MEM[20096];
assign MEM[28234] = MEM[19987] + MEM[20412];
assign MEM[28235] = MEM[19992] + MEM[20109];
assign MEM[28236] = MEM[19996] + MEM[20002];
assign MEM[28237] = MEM[19999] + MEM[20038];
assign MEM[28238] = MEM[20003] + MEM[20431];
assign MEM[28239] = MEM[20005] + MEM[20662];
assign MEM[28240] = MEM[20007] + MEM[20676];
assign MEM[28241] = MEM[20010] + MEM[20299];
assign MEM[28242] = MEM[20012] + MEM[20251];
assign MEM[28243] = MEM[20016] + MEM[20164];
assign MEM[28244] = MEM[20022] + MEM[20211];
assign MEM[28245] = MEM[20024] + MEM[20269];
assign MEM[28246] = MEM[20025] + MEM[20113];
assign MEM[28247] = MEM[20026] + MEM[20084];
assign MEM[28248] = MEM[20027] + MEM[20484];
assign MEM[28249] = MEM[20028] + MEM[20408];
assign MEM[28250] = MEM[20030] + MEM[20254];
assign MEM[28251] = MEM[20031] + MEM[21006];
assign MEM[28252] = MEM[20039] + MEM[20073];
assign MEM[28253] = MEM[20042] + MEM[20241];
assign MEM[28254] = MEM[20043] + MEM[20513];
assign MEM[28255] = MEM[20048] + MEM[20731];
assign MEM[28256] = MEM[20053] + MEM[20272];
assign MEM[28257] = MEM[20060] + MEM[20230];
assign MEM[28258] = MEM[20065] + MEM[20440];
assign MEM[28259] = MEM[20067] + MEM[20492];
assign MEM[28260] = MEM[20068] + MEM[20877];
assign MEM[28261] = MEM[20071] + MEM[20429];
assign MEM[28262] = MEM[20072] + MEM[20369];
assign MEM[28263] = MEM[20074] + MEM[20451];
assign MEM[28264] = MEM[20075] + MEM[20977];
assign MEM[28265] = MEM[20076] + MEM[20381];
assign MEM[28266] = MEM[20077] + MEM[20543];
assign MEM[28267] = MEM[20079] + MEM[20171];
assign MEM[28268] = MEM[20080] + MEM[20319];
assign MEM[28269] = MEM[20082] + MEM[20135];
assign MEM[28270] = MEM[20088] + MEM[20097];
assign MEM[28271] = MEM[20089] + MEM[21198];
assign MEM[28272] = MEM[20091] + MEM[20156];
assign MEM[28273] = MEM[20093] + MEM[20398];
assign MEM[28274] = MEM[20095] + MEM[20389];
assign MEM[28275] = MEM[20098] + MEM[20869];
assign MEM[28276] = MEM[20099] + MEM[20727];
assign MEM[28277] = MEM[20102] + MEM[20340];
assign MEM[28278] = MEM[20105] + MEM[20279];
assign MEM[28279] = MEM[20110] + MEM[20507];
assign MEM[28280] = MEM[20112] + MEM[20352];
assign MEM[28281] = MEM[20115] + MEM[20385];
assign MEM[28282] = MEM[20116] + MEM[20906];
assign MEM[28283] = MEM[20120] + MEM[20405];
assign MEM[28284] = MEM[20123] + MEM[20139];
assign MEM[28285] = MEM[20124] + MEM[20470];
assign MEM[28286] = MEM[20125] + MEM[21064];
assign MEM[28287] = MEM[20126] + MEM[21068];
assign MEM[28288] = MEM[20127] + MEM[20226];
assign MEM[28289] = MEM[20132] + MEM[20260];
assign MEM[28290] = MEM[20133] + MEM[20392];
assign MEM[28291] = MEM[20134] + MEM[20262];
assign MEM[28292] = MEM[20143] + MEM[20638];
assign MEM[28293] = MEM[20144] + MEM[20500];
assign MEM[28294] = MEM[20146] + MEM[20849];
assign MEM[28295] = MEM[20148] + MEM[20166];
assign MEM[28296] = MEM[20149] + MEM[21646];
assign MEM[28297] = MEM[20151] + MEM[20318];
assign MEM[28298] = MEM[20153] + MEM[20512];
assign MEM[28299] = MEM[20154] + MEM[20227];
assign MEM[28300] = MEM[20155] + MEM[20232];
assign MEM[28301] = MEM[20157] + MEM[20407];
assign MEM[28302] = MEM[20158] + MEM[20298];
assign MEM[28303] = MEM[20159] + MEM[20332];
assign MEM[28304] = MEM[20162] + MEM[20437];
assign MEM[28305] = MEM[20165] + MEM[20499];
assign MEM[28306] = MEM[20170] + MEM[20193];
assign MEM[28307] = MEM[20172] + MEM[20173];
assign MEM[28308] = MEM[20174] + MEM[20728];
assign MEM[28309] = MEM[20175] + MEM[20438];
assign MEM[28310] = MEM[20177] + MEM[20459];
assign MEM[28311] = MEM[20181] + MEM[20605];
assign MEM[28312] = MEM[20183] + MEM[20712];
assign MEM[28313] = MEM[20184] + MEM[20415];
assign MEM[28314] = MEM[20187] + MEM[20487];
assign MEM[28315] = MEM[20188] + MEM[20330];
assign MEM[28316] = MEM[20192] + MEM[20629];
assign MEM[28317] = MEM[20194] + MEM[21333];
assign MEM[28318] = MEM[20195] + MEM[20692];
assign MEM[28319] = MEM[20196] + MEM[21029];
assign MEM[28320] = MEM[20199] + MEM[20413];
assign MEM[28321] = MEM[20201] + MEM[20229];
assign MEM[28322] = MEM[20205] + MEM[20444];
assign MEM[28323] = MEM[20206] + MEM[20959];
assign MEM[28324] = MEM[20207] + MEM[20295];
assign MEM[28325] = MEM[20209] + MEM[20450];
assign MEM[28326] = MEM[20210] + MEM[20469];
assign MEM[28327] = MEM[20212] + MEM[20316];
assign MEM[28328] = MEM[20213] + MEM[20380];
assign MEM[28329] = MEM[20214] + MEM[20608];
assign MEM[28330] = MEM[20216] + MEM[20246];
assign MEM[28331] = MEM[20217] + MEM[20224];
assign MEM[28332] = MEM[20219] + MEM[20715];
assign MEM[28333] = MEM[20220] + MEM[20321];
assign MEM[28334] = MEM[20228] + MEM[20338];
assign MEM[28335] = MEM[20231] + MEM[20243];
assign MEM[28336] = MEM[20233] + MEM[20571];
assign MEM[28337] = MEM[20234] + MEM[20326];
assign MEM[28338] = MEM[20237] + MEM[20962];
assign MEM[28339] = MEM[20238] + MEM[20515];
assign MEM[28340] = MEM[20239] + MEM[20436];
assign MEM[28341] = MEM[20248] + MEM[20305];
assign MEM[28342] = MEM[20249] + MEM[20522];
assign MEM[28343] = MEM[20250] + MEM[20458];
assign MEM[28344] = MEM[20257] + MEM[20573];
assign MEM[28345] = MEM[20261] + MEM[20466];
assign MEM[28346] = MEM[20263] + MEM[20675];
assign MEM[28347] = MEM[20264] + MEM[20418];
assign MEM[28348] = MEM[20267] + MEM[20327];
assign MEM[28349] = MEM[20275] + MEM[21301];
assign MEM[28350] = MEM[20276] + MEM[20823];
assign MEM[28351] = MEM[20277] + MEM[20403];
assign MEM[28352] = MEM[20281] + MEM[20375];
assign MEM[28353] = MEM[20285] + MEM[21075];
assign MEM[28354] = MEM[20288] + MEM[20336];
assign MEM[28355] = MEM[20289] + MEM[21741];
assign MEM[28356] = MEM[20290] + MEM[20296];
assign MEM[28357] = MEM[20292] + MEM[20475];
assign MEM[28358] = MEM[20293] + MEM[20333];
assign MEM[28359] = MEM[20302] + MEM[21084];
assign MEM[28360] = MEM[20303] + MEM[20616];
assign MEM[28361] = MEM[20306] + MEM[20434];
assign MEM[28362] = MEM[20307] + MEM[20442];
assign MEM[28363] = MEM[20308] + MEM[20942];
assign MEM[28364] = MEM[20309] + MEM[20528];
assign MEM[28365] = MEM[20310] + MEM[20311];
assign MEM[28366] = MEM[20313] + MEM[20866];
assign MEM[28367] = MEM[20315] + MEM[20324];
assign MEM[28368] = MEM[20317] + MEM[20599];
assign MEM[28369] = MEM[20320] + MEM[20987];
assign MEM[28370] = MEM[20322] + MEM[20627];
assign MEM[28371] = MEM[20323] + MEM[20619];
assign MEM[28372] = MEM[20328] + MEM[20567];
assign MEM[28373] = MEM[20331] + MEM[20659];
assign MEM[28374] = MEM[20334] + MEM[20597];
assign MEM[28375] = MEM[20335] + MEM[20773];
assign MEM[28376] = MEM[20337] + MEM[20545];
assign MEM[28377] = MEM[20339] + MEM[21211];
assign MEM[28378] = MEM[20341] + MEM[20468];
assign MEM[28379] = MEM[20343] + MEM[20596];
assign MEM[28380] = MEM[20344] + MEM[21158];
assign MEM[28381] = MEM[20346] + MEM[20556];
assign MEM[28382] = MEM[20347] + MEM[20503];
assign MEM[28383] = MEM[20353] + MEM[20630];
assign MEM[28384] = MEM[20354] + MEM[20610];
assign MEM[28385] = MEM[20356] + MEM[20695];
assign MEM[28386] = MEM[20357] + MEM[20606];
assign MEM[28387] = MEM[20358] + MEM[20461];
assign MEM[28388] = MEM[20359] + MEM[20361];
assign MEM[28389] = MEM[20360] + MEM[20617];
assign MEM[28390] = MEM[20364] + MEM[20551];
assign MEM[28391] = MEM[20365] + MEM[20497];
assign MEM[28392] = MEM[20367] + MEM[20410];
assign MEM[28393] = MEM[20370] + MEM[21338];
assign MEM[28394] = MEM[20371] + MEM[20800];
assign MEM[28395] = MEM[20377] + MEM[20579];
assign MEM[28396] = MEM[20379] + MEM[20755];
assign MEM[28397] = MEM[20382] + MEM[20406];
assign MEM[28398] = MEM[20383] + MEM[20553];
assign MEM[28399] = MEM[20388] + MEM[20552];
assign MEM[28400] = MEM[20390] + MEM[21023];
assign MEM[28401] = MEM[20391] + MEM[20741];
assign MEM[28402] = MEM[20393] + MEM[20397];
assign MEM[28403] = MEM[20395] + MEM[20448];
assign MEM[28404] = MEM[20396] + MEM[20813];
assign MEM[28405] = MEM[20401] + MEM[20669];
assign MEM[28406] = MEM[20402] + MEM[20956];
assign MEM[28407] = MEM[20404] + MEM[20625];
assign MEM[28408] = MEM[20411] + MEM[20524];
assign MEM[28409] = MEM[20416] + MEM[21079];
assign MEM[28410] = MEM[20417] + MEM[20430];
assign MEM[28411] = MEM[20419] + MEM[20566];
assign MEM[28412] = MEM[20423] + MEM[20691];
assign MEM[28413] = MEM[20424] + MEM[20753];
assign MEM[28414] = MEM[20425] + MEM[20804];
assign MEM[28415] = MEM[20432] + MEM[21116];
assign MEM[28416] = MEM[20435] + MEM[20439];
assign MEM[28417] = MEM[20443] + MEM[20501];
assign MEM[28418] = MEM[20445] + MEM[20637];
assign MEM[28419] = MEM[20449] + MEM[20688];
assign MEM[28420] = MEM[20452] + MEM[21154];
assign MEM[28421] = MEM[20453] + MEM[20639];
assign MEM[28422] = MEM[20454] + MEM[20534];
assign MEM[28423] = MEM[20456] + MEM[21351];
assign MEM[28424] = MEM[20464] + MEM[22059];
assign MEM[28425] = MEM[20465] + MEM[20995];
assign MEM[28426] = MEM[20467] + MEM[21282];
assign MEM[28427] = MEM[20471] + MEM[21004];
assign MEM[28428] = MEM[20472] + MEM[20793];
assign MEM[28429] = MEM[20482] + MEM[21054];
assign MEM[28430] = MEM[20483] + MEM[20641];
assign MEM[28431] = MEM[20485] + MEM[20634];
assign MEM[28432] = MEM[20488] + MEM[20520];
assign MEM[28433] = MEM[20489] + MEM[20725];
assign MEM[28434] = MEM[20498] + MEM[21132];
assign MEM[28435] = MEM[20502] + MEM[20873];
assign MEM[28436] = MEM[20504] + MEM[20928];
assign MEM[28437] = MEM[20505] + MEM[21448];
assign MEM[28438] = MEM[20506] + MEM[20665];
assign MEM[28439] = MEM[20509] + MEM[20594];
assign MEM[28440] = MEM[20510] + MEM[21049];
assign MEM[28441] = MEM[20511] + MEM[20590];
assign MEM[28442] = MEM[20517] + MEM[21220];
assign MEM[28443] = MEM[20518] + MEM[21051];
assign MEM[28444] = MEM[20519] + MEM[20796];
assign MEM[28445] = MEM[20525] + MEM[20818];
assign MEM[28446] = MEM[20526] + MEM[20541];
assign MEM[28447] = MEM[20527] + MEM[20834];
assign MEM[28448] = MEM[20529] + MEM[20709];
assign MEM[28449] = MEM[20530] + MEM[20925];
assign MEM[28450] = MEM[20531] + MEM[20948];
assign MEM[28451] = MEM[20533] + MEM[21753];
assign MEM[28452] = MEM[20537] + MEM[20859];
assign MEM[28453] = MEM[20538] + MEM[20626];
assign MEM[28454] = MEM[20542] + MEM[20726];
assign MEM[28455] = MEM[20544] + MEM[20756];
assign MEM[28456] = MEM[20546] + MEM[20843];
assign MEM[28457] = MEM[20548] + MEM[20585];
assign MEM[28458] = MEM[20549] + MEM[20583];
assign MEM[28459] = MEM[20554] + MEM[21072];
assign MEM[28460] = MEM[20555] + MEM[20704];
assign MEM[28461] = MEM[20560] + MEM[20887];
assign MEM[28462] = MEM[20562] + MEM[20730];
assign MEM[28463] = MEM[20563] + MEM[20654];
assign MEM[28464] = MEM[20565] + MEM[20774];
assign MEM[28465] = MEM[20568] + MEM[20680];
assign MEM[28466] = MEM[20570] + MEM[20612];
assign MEM[28467] = MEM[20572] + MEM[21159];
assign MEM[28468] = MEM[20574] + MEM[21234];
assign MEM[28469] = MEM[20576] + MEM[20799];
assign MEM[28470] = MEM[20577] + MEM[20926];
assign MEM[28471] = MEM[20578] + MEM[20600];
assign MEM[28472] = MEM[20580] + MEM[20614];
assign MEM[28473] = MEM[20581] + MEM[21200];
assign MEM[28474] = MEM[20582] + MEM[20848];
assign MEM[28475] = MEM[20586] + MEM[20896];
assign MEM[28476] = MEM[20587] + MEM[20722];
assign MEM[28477] = MEM[20588] + MEM[20952];
assign MEM[28478] = MEM[20591] + MEM[20672];
assign MEM[28479] = MEM[20593] + MEM[20777];
assign MEM[28480] = MEM[20595] + MEM[21467];
assign MEM[28481] = MEM[20601] + MEM[21092];
assign MEM[28482] = MEM[20603] + MEM[21390];
assign MEM[28483] = MEM[20604] + MEM[20808];
assign MEM[28484] = MEM[20607] + MEM[20862];
assign MEM[28485] = MEM[20613] + MEM[20618];
assign MEM[28486] = MEM[20615] + MEM[21574];
assign MEM[28487] = MEM[20620] + MEM[20652];
assign MEM[28488] = MEM[20621] + MEM[21292];
assign MEM[28489] = MEM[20624] + MEM[20826];
assign MEM[28490] = MEM[20628] + MEM[20658];
assign MEM[28491] = MEM[20631] + MEM[20679];
assign MEM[28492] = MEM[20633] + MEM[20841];
assign MEM[28493] = MEM[20636] + MEM[20650];
assign MEM[28494] = MEM[20642] + MEM[20713];
assign MEM[28495] = MEM[20643] + MEM[20807];
assign MEM[28496] = MEM[20644] + MEM[20754];
assign MEM[28497] = MEM[20645] + MEM[21454];
assign MEM[28498] = MEM[20646] + MEM[20931];
assign MEM[28499] = MEM[20647] + MEM[20747];
assign MEM[28500] = MEM[20648] + MEM[20982];
assign MEM[28501] = MEM[20651] + MEM[20949];
assign MEM[28502] = MEM[20653] + MEM[20683];
assign MEM[28503] = MEM[20655] + MEM[21133];
assign MEM[28504] = MEM[20656] + MEM[20868];
assign MEM[28505] = MEM[20660] + MEM[21314];
assign MEM[28506] = MEM[20663] + MEM[20790];
assign MEM[28507] = MEM[20666] + MEM[21238];
assign MEM[28508] = MEM[20667] + MEM[21318];
assign MEM[28509] = MEM[20668] + MEM[21131];
assign MEM[28510] = MEM[20670] + MEM[20945];
assign MEM[28511] = MEM[20674] + MEM[20707];
assign MEM[28512] = MEM[20677] + MEM[20888];
assign MEM[28513] = MEM[20678] + MEM[20861];
assign MEM[28514] = MEM[20684] + MEM[20708];
assign MEM[28515] = MEM[20685] + MEM[20851];
assign MEM[28516] = MEM[20686] + MEM[21178];
assign MEM[28517] = MEM[20687] + MEM[21192];
assign MEM[28518] = MEM[20689] + MEM[21328];
assign MEM[28519] = MEM[20690] + MEM[21446];
assign MEM[28520] = MEM[20698] + MEM[20802];
assign MEM[28521] = MEM[20700] + MEM[20855];
assign MEM[28522] = MEM[20702] + MEM[20738];
assign MEM[28523] = MEM[20705] + MEM[20806];
assign MEM[28524] = MEM[20710] + MEM[20746];
assign MEM[28525] = MEM[20711] + MEM[21562];
assign MEM[28526] = MEM[20717] + MEM[20935];
assign MEM[28527] = MEM[20718] + MEM[20763];
assign MEM[28528] = MEM[20719] + MEM[20760];
assign MEM[28529] = MEM[20720] + MEM[20788];
assign MEM[28530] = MEM[20721] + MEM[21756];
assign MEM[28531] = MEM[20723] + MEM[21048];
assign MEM[28532] = MEM[20724] + MEM[20776];
assign MEM[28533] = MEM[20729] + MEM[21129];
assign MEM[28534] = MEM[20732] + MEM[21036];
assign MEM[28535] = MEM[20733] + MEM[21488];
assign MEM[28536] = MEM[20734] + MEM[20903];
assign MEM[28537] = MEM[20735] + MEM[20828];
assign MEM[28538] = MEM[20736] + MEM[20783];
assign MEM[28539] = MEM[20739] + MEM[20805];
assign MEM[28540] = MEM[20743] + MEM[20779];
assign MEM[28541] = MEM[20744] + MEM[21355];
assign MEM[28542] = MEM[20745] + MEM[21089];
assign MEM[28543] = MEM[20748] + MEM[20852];
assign MEM[28544] = MEM[20750] + MEM[20915];
assign MEM[28545] = MEM[20751] + MEM[20798];
assign MEM[28546] = MEM[20758] + MEM[21153];
assign MEM[28547] = MEM[20759] + MEM[20976];
assign MEM[28548] = MEM[20762] + MEM[20803];
assign MEM[28549] = MEM[20766] + MEM[21106];
assign MEM[28550] = MEM[20767] + MEM[20801];
assign MEM[28551] = MEM[20771] + MEM[21056];
assign MEM[28552] = MEM[20778] + MEM[21014];
assign MEM[28553] = MEM[20781] + MEM[21169];
assign MEM[28554] = MEM[20787] + MEM[21261];
assign MEM[28555] = MEM[20789] + MEM[21052];
assign MEM[28556] = MEM[20791] + MEM[20810];
assign MEM[28557] = MEM[20792] + MEM[21176];
assign MEM[28558] = MEM[20794] + MEM[20836];
assign MEM[28559] = MEM[20797] + MEM[21786];
assign MEM[28560] = MEM[20809] + MEM[20833];
assign MEM[28561] = MEM[20811] + MEM[21286];
assign MEM[28562] = MEM[20814] + MEM[20996];
assign MEM[28563] = MEM[20816] + MEM[21081];
assign MEM[28564] = MEM[20819] + MEM[21298];
assign MEM[28565] = MEM[20820] + MEM[20824];
assign MEM[28566] = MEM[20822] + MEM[20932];
assign MEM[28567] = MEM[20825] + MEM[21168];
assign MEM[28568] = MEM[20827] + MEM[20898];
assign MEM[28569] = MEM[20829] + MEM[21358];
assign MEM[28570] = MEM[20830] + MEM[20883];
assign MEM[28571] = MEM[20832] + MEM[20966];
assign MEM[28572] = MEM[20835] + MEM[21204];
assign MEM[28573] = MEM[20837] + MEM[21223];
assign MEM[28574] = MEM[20838] + MEM[20894];
assign MEM[28575] = MEM[20839] + MEM[21680];
assign MEM[28576] = MEM[20840] + MEM[21660];
assign MEM[28577] = MEM[20842] + MEM[20882];
assign MEM[28578] = MEM[20844] + MEM[21101];
assign MEM[28579] = MEM[20850] + MEM[21942];
assign MEM[28580] = MEM[20853] + MEM[21697];
assign MEM[28581] = MEM[20854] + MEM[21174];
assign MEM[28582] = MEM[20856] + MEM[21486];
assign MEM[28583] = MEM[20864] + MEM[21207];
assign MEM[28584] = MEM[20865] + MEM[21011];
assign MEM[28585] = MEM[20867] + MEM[21152];
assign MEM[28586] = MEM[20870] + MEM[21137];
assign MEM[28587] = MEM[20871] + MEM[21678];
assign MEM[28588] = MEM[20872] + MEM[21016];
assign MEM[28589] = MEM[20874] + MEM[20985];
assign MEM[28590] = MEM[20875] + MEM[21509];
assign MEM[28591] = MEM[20876] + MEM[21025];
assign MEM[28592] = MEM[20878] + MEM[20922];
assign MEM[28593] = MEM[20879] + MEM[20968];
assign MEM[28594] = MEM[20881] + MEM[21109];
assign MEM[28595] = MEM[20884] + MEM[20900];
assign MEM[28596] = MEM[20885] + MEM[20938];
assign MEM[28597] = MEM[20886] + MEM[20960];
assign MEM[28598] = MEM[20889] + MEM[21028];
assign MEM[28599] = MEM[20891] + MEM[21053];
assign MEM[28600] = MEM[20892] + MEM[21539];
assign MEM[28601] = MEM[20895] + MEM[21359];
assign MEM[28602] = MEM[20897] + MEM[21009];
assign MEM[28603] = MEM[20901] + MEM[21310];
assign MEM[28604] = MEM[20902] + MEM[20964];
assign MEM[28605] = MEM[20905] + MEM[21368];
assign MEM[28606] = MEM[20907] + MEM[21892];
assign MEM[28607] = MEM[20908] + MEM[21085];
assign MEM[28608] = MEM[20909] + MEM[21396];
assign MEM[28609] = MEM[20910] + MEM[21065];
assign MEM[28610] = MEM[20911] + MEM[21003];
assign MEM[28611] = MEM[20912] + MEM[21489];
assign MEM[28612] = MEM[20913] + MEM[21097];
assign MEM[28613] = MEM[20917] + MEM[21111];
assign MEM[28614] = MEM[20918] + MEM[21508];
assign MEM[28615] = MEM[20920] + MEM[21194];
assign MEM[28616] = MEM[20924] + MEM[21531];
assign MEM[28617] = MEM[20927] + MEM[20991];
assign MEM[28618] = MEM[20929] + MEM[20992];
assign MEM[28619] = MEM[20934] + MEM[20941];
assign MEM[28620] = MEM[20936] + MEM[21477];
assign MEM[28621] = MEM[20939] + MEM[21039];
assign MEM[28622] = MEM[20940] + MEM[21042];
assign MEM[28623] = MEM[20943] + MEM[21189];
assign MEM[28624] = MEM[20946] + MEM[21284];
assign MEM[28625] = MEM[20947] + MEM[21346];
assign MEM[28626] = MEM[20950] + MEM[21190];
assign MEM[28627] = MEM[20951] + MEM[21201];
assign MEM[28628] = MEM[20953] + MEM[21402];
assign MEM[28629] = MEM[20957] + MEM[21290];
assign MEM[28630] = MEM[20958] + MEM[21059];
assign MEM[28631] = MEM[20961] + MEM[21589];
assign MEM[28632] = MEM[20963] + MEM[21299];
assign MEM[28633] = MEM[20967] + MEM[21754];
assign MEM[28634] = MEM[20969] + MEM[21196];
assign MEM[28635] = MEM[20970] + MEM[21205];
assign MEM[28636] = MEM[20971] + MEM[21932];
assign MEM[28637] = MEM[20972] + MEM[21672];
assign MEM[28638] = MEM[20973] + MEM[21230];
assign MEM[28639] = MEM[20975] + MEM[22009];
assign MEM[28640] = MEM[20978] + MEM[21163];
assign MEM[28641] = MEM[20979] + MEM[21144];
assign MEM[28642] = MEM[20980] + MEM[21316];
assign MEM[28643] = MEM[20981] + MEM[21105];
assign MEM[28644] = MEM[20983] + MEM[21360];
assign MEM[28645] = MEM[20984] + MEM[21138];
assign MEM[28646] = MEM[20986] + MEM[21215];
assign MEM[28647] = MEM[20989] + MEM[21393];
assign MEM[28648] = MEM[20990] + MEM[21216];
assign MEM[28649] = MEM[20993] + MEM[21656];
assign MEM[28650] = MEM[20994] + MEM[21134];
assign MEM[28651] = MEM[20997] + MEM[21983];
assign MEM[28652] = MEM[20998] + MEM[21050];
assign MEM[28653] = MEM[20999] + MEM[21120];
assign MEM[28654] = MEM[21000] + MEM[21162];
assign MEM[28655] = MEM[21001] + MEM[21623];
assign MEM[28656] = MEM[21002] + MEM[21621];
assign MEM[28657] = MEM[21005] + MEM[21074];
assign MEM[28658] = MEM[21008] + MEM[21043];
assign MEM[28659] = MEM[21010] + MEM[21452];
assign MEM[28660] = MEM[21012] + MEM[21161];
assign MEM[28661] = MEM[21013] + MEM[21493];
assign MEM[28662] = MEM[21015] + MEM[21171];
assign MEM[28663] = MEM[21017] + MEM[21458];
assign MEM[28664] = MEM[21018] + MEM[21387];
assign MEM[28665] = MEM[21019] + MEM[21321];
assign MEM[28666] = MEM[21020] + MEM[21119];
assign MEM[28667] = MEM[21021] + MEM[21339];
assign MEM[28668] = MEM[21022] + MEM[21115];
assign MEM[28669] = MEM[21024] + MEM[21122];
assign MEM[28670] = MEM[21030] + MEM[21350];
assign MEM[28671] = MEM[21031] + MEM[21565];
assign MEM[28672] = MEM[21032] + MEM[21408];
assign MEM[28673] = MEM[21033] + MEM[21035];
assign MEM[28674] = MEM[21034] + MEM[21288];
assign MEM[28675] = MEM[21038] + MEM[21828];
assign MEM[28676] = MEM[21040] + MEM[21383];
assign MEM[28677] = MEM[21041] + MEM[21326];
assign MEM[28678] = MEM[21044] + MEM[21309];
assign MEM[28679] = MEM[21045] + MEM[21497];
assign MEM[28680] = MEM[21046] + MEM[21102];
assign MEM[28681] = MEM[21047] + MEM[21148];
assign MEM[28682] = MEM[21057] + MEM[21252];
assign MEM[28683] = MEM[21060] + MEM[21128];
assign MEM[28684] = MEM[21062] + MEM[21500];
assign MEM[28685] = MEM[21063] + MEM[21240];
assign MEM[28686] = MEM[21069] + MEM[21151];
assign MEM[28687] = MEM[21071] + MEM[21638];
assign MEM[28688] = MEM[21073] + MEM[21523];
assign MEM[28689] = MEM[21077] + MEM[21572];
assign MEM[28690] = MEM[21078] + MEM[21183];
assign MEM[28691] = MEM[21080] + MEM[21247];
assign MEM[28692] = MEM[21083] + MEM[21334];
assign MEM[28693] = MEM[21086] + MEM[22339];
assign MEM[28694] = MEM[21087] + MEM[21274];
assign MEM[28695] = MEM[21088] + MEM[21209];
assign MEM[28696] = MEM[21090] + MEM[21214];
assign MEM[28697] = MEM[21093] + MEM[21599];
assign MEM[28698] = MEM[21094] + MEM[21142];
assign MEM[28699] = MEM[21098] + MEM[21306];
assign MEM[28700] = MEM[21099] + MEM[21130];
assign MEM[28701] = MEM[21112] + MEM[21401];
assign MEM[28702] = MEM[21113] + MEM[21370];
assign MEM[28703] = MEM[21117] + MEM[21373];
assign MEM[28704] = MEM[21118] + MEM[21625];
assign MEM[28705] = MEM[21123] + MEM[21199];
assign MEM[28706] = MEM[21124] + MEM[21421];
assign MEM[28707] = MEM[21125] + MEM[21335];
assign MEM[28708] = MEM[21126] + MEM[21241];
assign MEM[28709] = MEM[21135] + MEM[21485];
assign MEM[28710] = MEM[21139] + MEM[21208];
assign MEM[28711] = MEM[21140] + MEM[21233];
assign MEM[28712] = MEM[21141] + MEM[21218];
assign MEM[28713] = MEM[21143] + MEM[21186];
assign MEM[28714] = MEM[21145] + MEM[21406];
assign MEM[28715] = MEM[21146] + MEM[21575];
assign MEM[28716] = MEM[21147] + MEM[21747];
assign MEM[28717] = MEM[21149] + MEM[21317];
assign MEM[28718] = MEM[21150] + MEM[21193];
assign MEM[28719] = MEM[21155] + MEM[21425];
assign MEM[28720] = MEM[21156] + MEM[21302];
assign MEM[28721] = MEM[21157] + MEM[21514];
assign MEM[28722] = MEM[21160] + MEM[21291];
assign MEM[28723] = MEM[21165] + MEM[21323];
assign MEM[28724] = MEM[21166] + MEM[21515];
assign MEM[28725] = MEM[21167] + MEM[21440];
assign MEM[28726] = MEM[21170] + MEM[21444];
assign MEM[28727] = MEM[21172] + MEM[21546];
assign MEM[28728] = MEM[21173] + MEM[21584];
assign MEM[28729] = MEM[21175] + MEM[21506];
assign MEM[28730] = MEM[21177] + MEM[21443];
assign MEM[28731] = MEM[21179] + MEM[21502];
assign MEM[28732] = MEM[21180] + MEM[21253];
assign MEM[28733] = MEM[21182] + MEM[21433];
assign MEM[28734] = MEM[21184] + MEM[21254];
assign MEM[28735] = MEM[21187] + MEM[21263];
assign MEM[28736] = MEM[21188] + MEM[21257];
assign MEM[28737] = MEM[21191] + MEM[21815];
assign MEM[28738] = MEM[21197] + MEM[22164];
assign MEM[28739] = MEM[21202] + MEM[21271];
assign MEM[28740] = MEM[21203] + MEM[21525];
assign MEM[28741] = MEM[21206] + MEM[21308];
assign MEM[28742] = MEM[21213] + MEM[21382];
assign MEM[28743] = MEM[21217] + MEM[21579];
assign MEM[28744] = MEM[21221] + MEM[21397];
assign MEM[28745] = MEM[21222] + MEM[21237];
assign MEM[28746] = MEM[21224] + MEM[21551];
assign MEM[28747] = MEM[21225] + MEM[21691];
assign MEM[28748] = MEM[21226] + MEM[21319];
assign MEM[28749] = MEM[21228] + MEM[21668];
assign MEM[28750] = MEM[21231] + MEM[21451];
assign MEM[28751] = MEM[21235] + MEM[21555];
assign MEM[28752] = MEM[21239] + MEM[21600];
assign MEM[28753] = MEM[21243] + MEM[21431];
assign MEM[28754] = MEM[21244] + MEM[21389];
assign MEM[28755] = MEM[21245] + MEM[21613];
assign MEM[28756] = MEM[21246] + MEM[21715];
assign MEM[28757] = MEM[21249] + MEM[21293];
assign MEM[28758] = MEM[21250] + MEM[21585];
assign MEM[28759] = MEM[21251] + MEM[21507];
assign MEM[28760] = MEM[21256] + MEM[21259];
assign MEM[28761] = MEM[21258] + MEM[21580];
assign MEM[28762] = MEM[21262] + MEM[21280];
assign MEM[28763] = MEM[21265] + MEM[21422];
assign MEM[28764] = MEM[21266] + MEM[21482];
assign MEM[28765] = MEM[21267] + MEM[21349];
assign MEM[28766] = MEM[21268] + MEM[22195];
assign MEM[28767] = MEM[21269] + MEM[22067];
assign MEM[28768] = MEM[21270] + MEM[21281];
assign MEM[28769] = MEM[21272] + MEM[21608];
assign MEM[28770] = MEM[21273] + MEM[21602];
assign MEM[28771] = MEM[21275] + MEM[21654];
assign MEM[28772] = MEM[21276] + MEM[22290];
assign MEM[28773] = MEM[21277] + MEM[21843];
assign MEM[28774] = MEM[21278] + MEM[21780];
assign MEM[28775] = MEM[21279] + MEM[21480];
assign MEM[28776] = MEM[21283] + MEM[21439];
assign MEM[28777] = MEM[21285] + MEM[22162];
assign MEM[28778] = MEM[21287] + MEM[22050];
assign MEM[28779] = MEM[21289] + MEM[21429];
assign MEM[28780] = MEM[21297] + MEM[21834];
assign MEM[28781] = MEM[21300] + MEM[21586];
assign MEM[28782] = MEM[21312] + MEM[21391];
assign MEM[28783] = MEM[21315] + MEM[21612];
assign MEM[28784] = MEM[21320] + MEM[21979];
assign MEM[28785] = MEM[21325] + MEM[21630];
assign MEM[28786] = MEM[21327] + MEM[21899];
assign MEM[28787] = MEM[21330] + MEM[21569];
assign MEM[28788] = MEM[21332] + MEM[21615];
assign MEM[28789] = MEM[21336] + MEM[21384];
assign MEM[28790] = MEM[21337] + MEM[21962];
assign MEM[28791] = MEM[21340] + MEM[21813];
assign MEM[28792] = MEM[21342] + MEM[21435];
assign MEM[28793] = MEM[21343] + MEM[22223];
assign MEM[28794] = MEM[21344] + MEM[21361];
assign MEM[28795] = MEM[21345] + MEM[21438];
assign MEM[28796] = MEM[21347] + MEM[21470];
assign MEM[28797] = MEM[21352] + MEM[21652];
assign MEM[28798] = MEM[21356] + MEM[21921];
assign MEM[28799] = MEM[21357] + MEM[22006];
assign MEM[28800] = MEM[21362] + MEM[21594];
assign MEM[28801] = MEM[21364] + MEM[21714];
assign MEM[28802] = MEM[21365] + MEM[21644];
assign MEM[28803] = MEM[21366] + MEM[22245];
assign MEM[28804] = MEM[21367] + MEM[21417];
assign MEM[28805] = MEM[21374] + MEM[21447];
assign MEM[28806] = MEM[21375] + MEM[21527];
assign MEM[28807] = MEM[21377] + MEM[21739];
assign MEM[28808] = MEM[21378] + MEM[22151];
assign MEM[28809] = MEM[21379] + MEM[21491];
assign MEM[28810] = MEM[21380] + MEM[21951];
assign MEM[28811] = MEM[21385] + MEM[21823];
assign MEM[28812] = MEM[21388] + MEM[21392];
assign MEM[28813] = MEM[21395] + MEM[21423];
assign MEM[28814] = MEM[21398] + MEM[21563];
assign MEM[28815] = MEM[21399] + MEM[22926];
assign MEM[28816] = MEM[21400] + MEM[21468];
assign MEM[28817] = MEM[21403] + MEM[21434];
assign MEM[28818] = MEM[21405] + MEM[21677];
assign MEM[28819] = MEM[21407] + MEM[21821];
assign MEM[28820] = MEM[21409] + MEM[21721];
assign MEM[28821] = MEM[21410] + MEM[21542];
assign MEM[28822] = MEM[21411] + MEM[22081];
assign MEM[28823] = MEM[21412] + MEM[21726];
assign MEM[28824] = MEM[21413] + MEM[21550];
assign MEM[28825] = MEM[21414] + MEM[21946];
assign MEM[28826] = MEM[21415] + MEM[21496];
assign MEM[28827] = MEM[21416] + MEM[22526];
assign MEM[28828] = MEM[21419] + MEM[21830];
assign MEM[28829] = MEM[21420] + MEM[21475];
assign MEM[28830] = MEM[21424] + MEM[21890];
assign MEM[28831] = MEM[21426] + MEM[21478];
assign MEM[28832] = MEM[21427] + MEM[21681];
assign MEM[28833] = MEM[21432] + MEM[21793];
assign MEM[28834] = MEM[21437] + MEM[21926];
assign MEM[28835] = MEM[21441] + MEM[22294];
assign MEM[28836] = MEM[21442] + MEM[21499];
assign MEM[28837] = MEM[21450] + MEM[21568];
assign MEM[28838] = MEM[21455] + MEM[21505];
assign MEM[28839] = MEM[21456] + MEM[21968];
assign MEM[28840] = MEM[21459] + MEM[21717];
assign MEM[28841] = MEM[21460] + MEM[21985];
assign MEM[28842] = MEM[21461] + MEM[21734];
assign MEM[28843] = MEM[21462] + MEM[22087];
assign MEM[28844] = MEM[21464] + MEM[21479];
assign MEM[28845] = MEM[21466] + MEM[21846];
assign MEM[28846] = MEM[21469] + MEM[21831];
assign MEM[28847] = MEM[21471] + MEM[22011];
assign MEM[28848] = MEM[21472] + MEM[21969];
assign MEM[28849] = MEM[21474] + MEM[21498];
assign MEM[28850] = MEM[21476] + MEM[21869];
assign MEM[28851] = MEM[21481] + MEM[21750];
assign MEM[28852] = MEM[21483] + MEM[21682];
assign MEM[28853] = MEM[21487] + MEM[21609];
assign MEM[28854] = MEM[21490] + MEM[21689];
assign MEM[28855] = MEM[21492] + MEM[21855];
assign MEM[28856] = MEM[21494] + MEM[21577];
assign MEM[28857] = MEM[21495] + MEM[21788];
assign MEM[28858] = MEM[21501] + MEM[21519];
assign MEM[28859] = MEM[21503] + MEM[21548];
assign MEM[28860] = MEM[21511] + MEM[21676];
assign MEM[28861] = MEM[21512] + MEM[21604];
assign MEM[28862] = MEM[21513] + MEM[21709];
assign MEM[28863] = MEM[21516] + MEM[21560];
assign MEM[28864] = MEM[21518] + MEM[21708];
assign MEM[28865] = MEM[21520] + MEM[21658];
assign MEM[28866] = MEM[21521] + MEM[21636];
assign MEM[28867] = MEM[21522] + MEM[21933];
assign MEM[28868] = MEM[21524] + MEM[22637];
assign MEM[28869] = MEM[21526] + MEM[21611];
assign MEM[28870] = MEM[21528] + MEM[21794];
assign MEM[28871] = MEM[21529] + MEM[21749];
assign MEM[28872] = MEM[21532] + MEM[21544];
assign MEM[28873] = MEM[21533] + MEM[22614];
assign MEM[28874] = MEM[21534] + MEM[21902];
assign MEM[28875] = MEM[21535] + MEM[21661];
assign MEM[28876] = MEM[21537] + MEM[21995];
assign MEM[28877] = MEM[21540] + MEM[21699];
assign MEM[28878] = MEM[21541] + MEM[21704];
assign MEM[28879] = MEM[21545] + MEM[21666];
assign MEM[28880] = MEM[21549] + MEM[21770];
assign MEM[28881] = MEM[21552] + MEM[21603];
assign MEM[28882] = MEM[21553] + MEM[22123];
assign MEM[28883] = MEM[21554] + MEM[21819];
assign MEM[28884] = MEM[21556] + MEM[21837];
assign MEM[28885] = MEM[21557] + MEM[21873];
assign MEM[28886] = MEM[21559] + MEM[21797];
assign MEM[28887] = MEM[21561] + MEM[21870];
assign MEM[28888] = MEM[21564] + MEM[21583];
assign MEM[28889] = MEM[21566] + MEM[22714];
assign MEM[28890] = MEM[21567] + MEM[22735];
assign MEM[28891] = MEM[21573] + MEM[21807];
assign MEM[28892] = MEM[21576] + MEM[22256];
assign MEM[28893] = MEM[21578] + MEM[21614];
assign MEM[28894] = MEM[21582] + MEM[22130];
assign MEM[28895] = MEM[21587] + MEM[21719];
assign MEM[28896] = MEM[21588] + MEM[22314];
assign MEM[28897] = MEM[21591] + MEM[21746];
assign MEM[28898] = MEM[21592] + MEM[21799];
assign MEM[28899] = MEM[21593] + MEM[22424];
assign MEM[28900] = MEM[21597] + MEM[21779];
assign MEM[28901] = MEM[21601] + MEM[21617];
assign MEM[28902] = MEM[21605] + MEM[21851];
assign MEM[28903] = MEM[21606] + MEM[21649];
assign MEM[28904] = MEM[21610] + MEM[21619];
assign MEM[28905] = MEM[21616] + MEM[21701];
assign MEM[28906] = MEM[21620] + MEM[21961];
assign MEM[28907] = MEM[21622] + MEM[21859];
assign MEM[28908] = MEM[21624] + MEM[21838];
assign MEM[28909] = MEM[21626] + MEM[21941];
assign MEM[28910] = MEM[21628] + MEM[21694];
assign MEM[28911] = MEM[21629] + MEM[21670];
assign MEM[28912] = MEM[21631] + MEM[21740];
assign MEM[28913] = MEM[21632] + MEM[21880];
assign MEM[28914] = MEM[21634] + MEM[21733];
assign MEM[28915] = MEM[21635] + MEM[21769];
assign MEM[28916] = MEM[21637] + MEM[22363];
assign MEM[28917] = MEM[21639] + MEM[21716];
assign MEM[28918] = MEM[21641] + MEM[21910];
assign MEM[28919] = MEM[21643] + MEM[21737];
assign MEM[28920] = MEM[21648] + MEM[21690];
assign MEM[28921] = MEM[21650] + MEM[21736];
assign MEM[28922] = MEM[21651] + MEM[21735];
assign MEM[28923] = MEM[21653] + MEM[21729];
assign MEM[28924] = MEM[21655] + MEM[21688];
assign MEM[28925] = MEM[21657] + MEM[21844];
assign MEM[28926] = MEM[21659] + MEM[21818];
assign MEM[28927] = MEM[21662] + MEM[21973];
assign MEM[28928] = MEM[21663] + MEM[21771];
assign MEM[28929] = MEM[21664] + MEM[21781];
assign MEM[28930] = MEM[21665] + MEM[22272];
assign MEM[28931] = MEM[21667] + MEM[23162];
assign MEM[28932] = MEM[21669] + MEM[22106];
assign MEM[28933] = MEM[21671] + MEM[21695];
assign MEM[28934] = MEM[21673] + MEM[21796];
assign MEM[28935] = MEM[21674] + MEM[21795];
assign MEM[28936] = MEM[21675] + MEM[21993];
assign MEM[28937] = MEM[21679] + MEM[21758];
assign MEM[28938] = MEM[21684] + MEM[21738];
assign MEM[28939] = MEM[21685] + MEM[21866];
assign MEM[28940] = MEM[21686] + MEM[21791];
assign MEM[28941] = MEM[21692] + MEM[22230];
assign MEM[28942] = MEM[21693] + MEM[22556];
assign MEM[28943] = MEM[21696] + MEM[21940];
assign MEM[28944] = MEM[21698] + MEM[21700];
assign MEM[28945] = MEM[21702] + MEM[21728];
assign MEM[28946] = MEM[21703] + MEM[22167];
assign MEM[28947] = MEM[21705] + MEM[21839];
assign MEM[28948] = MEM[21706] + MEM[22134];
assign MEM[28949] = MEM[21707] + MEM[22046];
assign MEM[28950] = MEM[21710] + MEM[21848];
assign MEM[28951] = MEM[21711] + MEM[21981];
assign MEM[28952] = MEM[21712] + MEM[21816];
assign MEM[28953] = MEM[21720] + MEM[21982];
assign MEM[28954] = MEM[21723] + MEM[21810];
assign MEM[28955] = MEM[21725] + MEM[22080];
assign MEM[28956] = MEM[21727] + MEM[21858];
assign MEM[28957] = MEM[21730] + MEM[22429];
assign MEM[28958] = MEM[21742] + MEM[22312];
assign MEM[28959] = MEM[21743] + MEM[22678];
assign MEM[28960] = MEM[21744] + MEM[21878];
assign MEM[28961] = MEM[21745] + MEM[22060];
assign MEM[28962] = MEM[21748] + MEM[21903];
assign MEM[28963] = MEM[21751] + MEM[21991];
assign MEM[28964] = MEM[21752] + MEM[21812];
assign MEM[28965] = MEM[21757] + MEM[21845];
assign MEM[28966] = MEM[21759] + MEM[21914];
assign MEM[28967] = MEM[21760] + MEM[22336];
assign MEM[28968] = MEM[21761] + MEM[21988];
assign MEM[28969] = MEM[21763] + MEM[22094];
assign MEM[28970] = MEM[21764] + MEM[22069];
assign MEM[28971] = MEM[21767] + MEM[22056];
assign MEM[28972] = MEM[21768] + MEM[21904];
assign MEM[28973] = MEM[21772] + MEM[22307];
assign MEM[28974] = MEM[21773] + MEM[22183];
assign MEM[28975] = MEM[21775] + MEM[22140];
assign MEM[28976] = MEM[21776] + MEM[21901];
assign MEM[28977] = MEM[21777] + MEM[22483];
assign MEM[28978] = MEM[21778] + MEM[21829];
assign MEM[28979] = MEM[21782] + MEM[21938];
assign MEM[28980] = MEM[21783] + MEM[22101];
assign MEM[28981] = MEM[21784] + MEM[22032];
assign MEM[28982] = MEM[21785] + MEM[22173];
assign MEM[28983] = MEM[21789] + MEM[22400];
assign MEM[28984] = MEM[21792] + MEM[21917];
assign MEM[28985] = MEM[21800] + MEM[21882];
assign MEM[28986] = MEM[21803] + MEM[21884];
assign MEM[28987] = MEM[21804] + MEM[22025];
assign MEM[28988] = MEM[21805] + MEM[22405];
assign MEM[28989] = MEM[21808] + MEM[21996];
assign MEM[28990] = MEM[21809] + MEM[22257];
assign MEM[28991] = MEM[21811] + MEM[22255];
assign MEM[28992] = MEM[21814] + MEM[21824];
assign MEM[28993] = MEM[21817] + MEM[21857];
assign MEM[28994] = MEM[21820] + MEM[21911];
assign MEM[28995] = MEM[21822] + MEM[22287];
assign MEM[28996] = MEM[21826] + MEM[21853];
assign MEM[28997] = MEM[21827] + MEM[21888];
assign MEM[28998] = MEM[21833] + MEM[22044];
assign MEM[28999] = MEM[21835] + MEM[21947];
assign MEM[29000] = MEM[21840] + MEM[22643];
assign MEM[29001] = MEM[21842] + MEM[22284];
assign MEM[29002] = MEM[21847] + MEM[22358];
assign MEM[29003] = MEM[21849] + MEM[22159];
assign MEM[29004] = MEM[21850] + MEM[22615];
assign MEM[29005] = MEM[21852] + MEM[22311];
assign MEM[29006] = MEM[21854] + MEM[22076];
assign MEM[29007] = MEM[21860] + MEM[22315];
assign MEM[29008] = MEM[21861] + MEM[22460];
assign MEM[29009] = MEM[21863] + MEM[22587];
assign MEM[29010] = MEM[21864] + MEM[22002];
assign MEM[29011] = MEM[21865] + MEM[22102];
assign MEM[29012] = MEM[21868] + MEM[21966];
assign MEM[29013] = MEM[21872] + MEM[22051];
assign MEM[29014] = MEM[21874] + MEM[22292];
assign MEM[29015] = MEM[21875] + MEM[22340];
assign MEM[29016] = MEM[21876] + MEM[22088];
assign MEM[29017] = MEM[21877] + MEM[21943];
assign MEM[29018] = MEM[21879] + MEM[22286];
assign MEM[29019] = MEM[21881] + MEM[22200];
assign MEM[29020] = MEM[21883] + MEM[22073];
assign MEM[29021] = MEM[21885] + MEM[22676];
assign MEM[29022] = MEM[21887] + MEM[21953];
assign MEM[29023] = MEM[21889] + MEM[22525];
assign MEM[29024] = MEM[21891] + MEM[22469];
assign MEM[29025] = MEM[21893] + MEM[22176];
assign MEM[29026] = MEM[21896] + MEM[21915];
assign MEM[29027] = MEM[21897] + MEM[21929];
assign MEM[29028] = MEM[21898] + MEM[22054];
assign MEM[29029] = MEM[21900] + MEM[22246];
assign MEM[29030] = MEM[21905] + MEM[22161];
assign MEM[29031] = MEM[21907] + MEM[22007];
assign MEM[29032] = MEM[21908] + MEM[22276];
assign MEM[29033] = MEM[21912] + MEM[22077];
assign MEM[29034] = MEM[21913] + MEM[21957];
assign MEM[29035] = MEM[21916] + MEM[21918];
assign MEM[29036] = MEM[21919] + MEM[22066];
assign MEM[29037] = MEM[21922] + MEM[22158];
assign MEM[29038] = MEM[21923] + MEM[22045];
assign MEM[29039] = MEM[21928] + MEM[22456];
assign MEM[29040] = MEM[21930] + MEM[22326];
assign MEM[29041] = MEM[21931] + MEM[22262];
assign MEM[29042] = MEM[21935] + MEM[21949];
assign MEM[29043] = MEM[21936] + MEM[22058];
assign MEM[29044] = MEM[21937] + MEM[22064];
assign MEM[29045] = MEM[21944] + MEM[22212];
assign MEM[29046] = MEM[21945] + MEM[22470];
assign MEM[29047] = MEM[21948] + MEM[22494];
assign MEM[29048] = MEM[21950] + MEM[22912];
assign MEM[29049] = MEM[21952] + MEM[22560];
assign MEM[29050] = MEM[21954] + MEM[22402];
assign MEM[29051] = MEM[21956] + MEM[22367];
assign MEM[29052] = MEM[21959] + MEM[22316];
assign MEM[29053] = MEM[21960] + MEM[22120];
assign MEM[29054] = MEM[21963] + MEM[22224];
assign MEM[29055] = MEM[21964] + MEM[22450];
assign MEM[29056] = MEM[21965] + MEM[22519];
assign MEM[29057] = MEM[21967] + MEM[22166];
assign MEM[29058] = MEM[21972] + MEM[22480];
assign MEM[29059] = MEM[21974] + MEM[22691];
assign MEM[29060] = MEM[21975] + MEM[22422];
assign MEM[29061] = MEM[21976] + MEM[22631];
assign MEM[29062] = MEM[21978] + MEM[22486];
assign MEM[29063] = MEM[21980] + MEM[21997];
assign MEM[29064] = MEM[21984] + MEM[22365];
assign MEM[29065] = MEM[21986] + MEM[22107];
assign MEM[29066] = MEM[21987] + MEM[22005];
assign MEM[29067] = MEM[21990] + MEM[22433];
assign MEM[29068] = MEM[21992] + MEM[22193];
assign MEM[29069] = MEM[21994] + MEM[22280];
assign MEM[29070] = MEM[21998] + MEM[23122];
assign MEM[29071] = MEM[21999] + MEM[22416];
assign MEM[29072] = MEM[22001] + MEM[22247];
assign MEM[29073] = MEM[22004] + MEM[22098];
assign MEM[29074] = MEM[22010] + MEM[22078];
assign MEM[29075] = MEM[22014] + MEM[22036];
assign MEM[29076] = MEM[22015] + MEM[22843];
assign MEM[29077] = MEM[22017] + MEM[22091];
assign MEM[29078] = MEM[22018] + MEM[22068];
assign MEM[29079] = MEM[22020] + MEM[22126];
assign MEM[29080] = MEM[22021] + MEM[23457];
assign MEM[29081] = MEM[22022] + MEM[22071];
assign MEM[29082] = MEM[22024] + MEM[22168];
assign MEM[29083] = MEM[22026] + MEM[22086];
assign MEM[29084] = MEM[22027] + MEM[22182];
assign MEM[29085] = MEM[22028] + MEM[22720];
assign MEM[29086] = MEM[22029] + MEM[22352];
assign MEM[29087] = MEM[22030] + MEM[22041];
assign MEM[29088] = MEM[22031] + MEM[22253];
assign MEM[29089] = MEM[22035] + MEM[22219];
assign MEM[29090] = MEM[22037] + MEM[22484];
assign MEM[29091] = MEM[22038] + MEM[22221];
assign MEM[29092] = MEM[22039] + MEM[22840];
assign MEM[29093] = MEM[22040] + MEM[22206];
assign MEM[29094] = MEM[22042] + MEM[22304];
assign MEM[29095] = MEM[22043] + MEM[23018];
assign MEM[29096] = MEM[22047] + MEM[22297];
assign MEM[29097] = MEM[22048] + MEM[22535];
assign MEM[29098] = MEM[22049] + MEM[22277];
assign MEM[29099] = MEM[22052] + MEM[22057];
assign MEM[29100] = MEM[22053] + MEM[22192];
assign MEM[29101] = MEM[22055] + MEM[22061];
assign MEM[29102] = MEM[22062] + MEM[22096];
assign MEM[29103] = MEM[22063] + MEM[22095];
assign MEM[29104] = MEM[22065] + MEM[22356];
assign MEM[29105] = MEM[22070] + MEM[22093];
assign MEM[29106] = MEM[22072] + MEM[22444];
assign MEM[29107] = MEM[22074] + MEM[22125];
assign MEM[29108] = MEM[22075] + MEM[22548];
assign MEM[29109] = MEM[22079] + MEM[22408];
assign MEM[29110] = MEM[22082] + MEM[22347];
assign MEM[29111] = MEM[22083] + MEM[22156];
assign MEM[29112] = MEM[22085] + MEM[22285];
assign MEM[29113] = MEM[22089] + MEM[22197];
assign MEM[29114] = MEM[22090] + MEM[22701];
assign MEM[29115] = MEM[22092] + MEM[22226];
assign MEM[29116] = MEM[22099] + MEM[22188];
assign MEM[29117] = MEM[22100] + MEM[22271];
assign MEM[29118] = MEM[22103] + MEM[22237];
assign MEM[29119] = MEM[22104] + MEM[22773];
assign MEM[29120] = MEM[22105] + MEM[22960];
assign MEM[29121] = MEM[22108] + MEM[22157];
assign MEM[29122] = MEM[22109] + MEM[22116];
assign MEM[29123] = MEM[22111] + MEM[22169];
assign MEM[29124] = MEM[22113] + MEM[22366];
assign MEM[29125] = MEM[22114] + MEM[22390];
assign MEM[29126] = MEM[22115] + MEM[22240];
assign MEM[29127] = MEM[22117] + MEM[22175];
assign MEM[29128] = MEM[22121] + MEM[22296];
assign MEM[29129] = MEM[22122] + MEM[24448];
assign MEM[29130] = MEM[22124] + MEM[22653];
assign MEM[29131] = MEM[22127] + MEM[22209];
assign MEM[29132] = MEM[22128] + MEM[22780];
assign MEM[29133] = MEM[22129] + MEM[22447];
assign MEM[29134] = MEM[22132] + MEM[22204];
assign MEM[29135] = MEM[22133] + MEM[22409];
assign MEM[29136] = MEM[22135] + MEM[22211];
assign MEM[29137] = MEM[22136] + MEM[22434];
assign MEM[29138] = MEM[22137] + MEM[22298];
assign MEM[29139] = MEM[22138] + MEM[22289];
assign MEM[29140] = MEM[22139] + MEM[22207];
assign MEM[29141] = MEM[22141] + MEM[22559];
assign MEM[29142] = MEM[22143] + MEM[22396];
assign MEM[29143] = MEM[22144] + MEM[22792];
assign MEM[29144] = MEM[22145] + MEM[22233];
assign MEM[29145] = MEM[22146] + MEM[22485];
assign MEM[29146] = MEM[22147] + MEM[22215];
assign MEM[29147] = MEM[22152] + MEM[24238];
assign MEM[29148] = MEM[22153] + MEM[22577];
assign MEM[29149] = MEM[22154] + MEM[23059];
assign MEM[29150] = MEM[22155] + MEM[23348];
assign MEM[29151] = MEM[22160] + MEM[22278];
assign MEM[29152] = MEM[22163] + MEM[22585];
assign MEM[29153] = MEM[22165] + MEM[22406];
assign MEM[29154] = MEM[22171] + MEM[22550];
assign MEM[29155] = MEM[22172] + MEM[22218];
assign MEM[29156] = MEM[22174] + MEM[22383];
assign MEM[29157] = MEM[22177] + MEM[22439];
assign MEM[29158] = MEM[22178] + MEM[22459];
assign MEM[29159] = MEM[22179] + MEM[22894];
assign MEM[29160] = MEM[22180] + MEM[22412];
assign MEM[29161] = MEM[22185] + MEM[22812];
assign MEM[29162] = MEM[22186] + MEM[22379];
assign MEM[29163] = MEM[22187] + MEM[22520];
assign MEM[29164] = MEM[22189] + MEM[22771];
assign MEM[29165] = MEM[22190] + MEM[23715];
assign MEM[29166] = MEM[22191] + MEM[22611];
assign MEM[29167] = MEM[22194] + MEM[22669];
assign MEM[29168] = MEM[22198] + MEM[22360];
assign MEM[29169] = MEM[22201] + MEM[22498];
assign MEM[29170] = MEM[22202] + MEM[22371];
assign MEM[29171] = MEM[22205] + MEM[22816];
assign MEM[29172] = MEM[22208] + MEM[22695];
assign MEM[29173] = MEM[22210] + MEM[22249];
assign MEM[29174] = MEM[22213] + MEM[22432];
assign MEM[29175] = MEM[22214] + MEM[22242];
assign MEM[29176] = MEM[22216] + MEM[22571];
assign MEM[29177] = MEM[22217] + MEM[22473];
assign MEM[29178] = MEM[22220] + MEM[22391];
assign MEM[29179] = MEM[22222] + MEM[22663];
assign MEM[29180] = MEM[22225] + MEM[22364];
assign MEM[29181] = MEM[22228] + MEM[23118];
assign MEM[29182] = MEM[22232] + MEM[22310];
assign MEM[29183] = MEM[22234] + MEM[22738];
assign MEM[29184] = MEM[22235] + MEM[22797];
assign MEM[29185] = MEM[22236] + MEM[22239];
assign MEM[29186] = MEM[22241] + MEM[22723];
assign MEM[29187] = MEM[22243] + MEM[22621];
assign MEM[29188] = MEM[22244] + MEM[22862];
assign MEM[29189] = MEM[22248] + MEM[22260];
assign MEM[29190] = MEM[22250] + MEM[22783];
assign MEM[29191] = MEM[22251] + MEM[23030];
assign MEM[29192] = MEM[22252] + MEM[22413];
assign MEM[29193] = MEM[22254] + MEM[22616];
assign MEM[29194] = MEM[22259] + MEM[22384];
assign MEM[29195] = MEM[22261] + MEM[22493];
assign MEM[29196] = MEM[22263] + MEM[22376];
assign MEM[29197] = MEM[22265] + MEM[22546];
assign MEM[29198] = MEM[22266] + MEM[22579];
assign MEM[29199] = MEM[22267] + MEM[22681];
assign MEM[29200] = MEM[22269] + MEM[22934];
assign MEM[29201] = MEM[22270] + MEM[23310];
assign MEM[29202] = MEM[22273] + MEM[22820];
assign MEM[29203] = MEM[22274] + MEM[22847];
assign MEM[29204] = MEM[22275] + MEM[22415];
assign MEM[29205] = MEM[22279] + MEM[22385];
assign MEM[29206] = MEM[22281] + MEM[22481];
assign MEM[29207] = MEM[22282] + MEM[22917];
assign MEM[29208] = MEM[22291] + MEM[22488];
assign MEM[29209] = MEM[22299] + MEM[22827];
assign MEM[29210] = MEM[22301] + MEM[22949];
assign MEM[29211] = MEM[22302] + MEM[22649];
assign MEM[29212] = MEM[22303] + MEM[22392];
assign MEM[29213] = MEM[22305] + MEM[22612];
assign MEM[29214] = MEM[22306] + MEM[22395];
assign MEM[29215] = MEM[22308] + MEM[22555];
assign MEM[29216] = MEM[22309] + MEM[22778];
assign MEM[29217] = MEM[22318] + MEM[22377];
assign MEM[29218] = MEM[22319] + MEM[22940];
assign MEM[29219] = MEM[22320] + MEM[22467];
assign MEM[29220] = MEM[22321] + MEM[22355];
assign MEM[29221] = MEM[22322] + MEM[22748];
assign MEM[29222] = MEM[22323] + MEM[22943];
assign MEM[29223] = MEM[22324] + MEM[22401];
assign MEM[29224] = MEM[22325] + MEM[22533];
assign MEM[29225] = MEM[22328] + MEM[22386];
assign MEM[29226] = MEM[22329] + MEM[23022];
assign MEM[29227] = MEM[22330] + MEM[22855];
assign MEM[29228] = MEM[22331] + MEM[23274];
assign MEM[29229] = MEM[22332] + MEM[22497];
assign MEM[29230] = MEM[22333] + MEM[22378];
assign MEM[29231] = MEM[22334] + MEM[22956];
assign MEM[29232] = MEM[22335] + MEM[23129];
assign MEM[29233] = MEM[22337] + MEM[22905];
assign MEM[29234] = MEM[22338] + MEM[22739];
assign MEM[29235] = MEM[22342] + MEM[22740];
assign MEM[29236] = MEM[22343] + MEM[22500];
assign MEM[29237] = MEM[22346] + MEM[22532];
assign MEM[29238] = MEM[22348] + MEM[22594];
assign MEM[29239] = MEM[22350] + MEM[22578];
assign MEM[29240] = MEM[22351] + MEM[23155];
assign MEM[29241] = MEM[22353] + MEM[22764];
assign MEM[29242] = MEM[22354] + MEM[22545];
assign MEM[29243] = MEM[22359] + MEM[22962];
assign MEM[29244] = MEM[22361] + MEM[23117];
assign MEM[29245] = MEM[22362] + MEM[22599];
assign MEM[29246] = MEM[22370] + MEM[22648];
assign MEM[29247] = MEM[22372] + MEM[22465];
assign MEM[29248] = MEM[22373] + MEM[22573];
assign MEM[29249] = MEM[22375] + MEM[22933];
assign MEM[29250] = MEM[22380] + MEM[22896];
assign MEM[29251] = MEM[22381] + MEM[22388];
assign MEM[29252] = MEM[22382] + MEM[22538];
assign MEM[29253] = MEM[22387] + MEM[22620];
assign MEM[29254] = MEM[22389] + MEM[22451];
assign MEM[29255] = MEM[22393] + MEM[22489];
assign MEM[29256] = MEM[22394] + MEM[22742];
assign MEM[29257] = MEM[22397] + MEM[22657];
assign MEM[29258] = MEM[22399] + MEM[22769];
assign MEM[29259] = MEM[22403] + MEM[23047];
assign MEM[29260] = MEM[22404] + MEM[22506];
assign MEM[29261] = MEM[22410] + MEM[22531];
assign MEM[29262] = MEM[22411] + MEM[22457];
assign MEM[29263] = MEM[22414] + MEM[22463];
assign MEM[29264] = MEM[22418] + MEM[22677];
assign MEM[29265] = MEM[22421] + MEM[22455];
assign MEM[29266] = MEM[22423] + MEM[23023];
assign MEM[29267] = MEM[22426] + MEM[22629];
assign MEM[29268] = MEM[22427] + MEM[24005];
assign MEM[29269] = MEM[22428] + MEM[22453];
assign MEM[29270] = MEM[22430] + MEM[22452];
assign MEM[29271] = MEM[22431] + MEM[22517];
assign MEM[29272] = MEM[22435] + MEM[22524];
assign MEM[29273] = MEM[22436] + MEM[22628];
assign MEM[29274] = MEM[22437] + MEM[22872];
assign MEM[29275] = MEM[22440] + MEM[22495];
assign MEM[29276] = MEM[22441] + MEM[22979];
assign MEM[29277] = MEM[22443] + MEM[22513];
assign MEM[29278] = MEM[22445] + MEM[22693];
assign MEM[29279] = MEM[22448] + MEM[22939];
assign MEM[29280] = MEM[22454] + MEM[22753];
assign MEM[29281] = MEM[22458] + MEM[22802];
assign MEM[29282] = MEM[22461] + MEM[22487];
assign MEM[29283] = MEM[22462] + MEM[22825];
assign MEM[29284] = MEM[22464] + MEM[23007];
assign MEM[29285] = MEM[22466] + MEM[22508];
assign MEM[29286] = MEM[22471] + MEM[22478];
assign MEM[29287] = MEM[22472] + MEM[22619];
assign MEM[29288] = MEM[22474] + MEM[22636];
assign MEM[29289] = MEM[22476] + MEM[23530];
assign MEM[29290] = MEM[22477] + MEM[22947];
assign MEM[29291] = MEM[22479] + MEM[22965];
assign MEM[29292] = MEM[22482] + MEM[23197];
assign MEM[29293] = MEM[22490] + MEM[23762];
assign MEM[29294] = MEM[22491] + MEM[22911];
assign MEM[29295] = MEM[22492] + MEM[22624];
assign MEM[29296] = MEM[22496] + MEM[22607];
assign MEM[29297] = MEM[22499] + MEM[22791];
assign MEM[29298] = MEM[22501] + MEM[23025];
assign MEM[29299] = MEM[22502] + MEM[22689];
assign MEM[29300] = MEM[22503] + MEM[22635];
assign MEM[29301] = MEM[22504] + MEM[22536];
assign MEM[29302] = MEM[22505] + MEM[22789];
assign MEM[29303] = MEM[22507] + MEM[22844];
assign MEM[29304] = MEM[22512] + MEM[23020];
assign MEM[29305] = MEM[22516] + MEM[22751];
assign MEM[29306] = MEM[22518] + MEM[22561];
assign MEM[29307] = MEM[22521] + MEM[22830];
assign MEM[29308] = MEM[22522] + MEM[22542];
assign MEM[29309] = MEM[22523] + MEM[22697];
assign MEM[29310] = MEM[22527] + MEM[22922];
assign MEM[29311] = MEM[22528] + MEM[22717];
assign MEM[29312] = MEM[22529] + MEM[22630];
assign MEM[29313] = MEM[22530] + MEM[22877];
assign MEM[29314] = MEM[22534] + MEM[22733];
assign MEM[29315] = MEM[22537] + MEM[22602];
assign MEM[29316] = MEM[22539] + MEM[22777];
assign MEM[29317] = MEM[22540] + MEM[22814];
assign MEM[29318] = MEM[22541] + MEM[22826];
assign MEM[29319] = MEM[22543] + MEM[22743];
assign MEM[29320] = MEM[22544] + MEM[22842];
assign MEM[29321] = MEM[22547] + MEM[23105];
assign MEM[29322] = MEM[22549] + MEM[22672];
assign MEM[29323] = MEM[22551] + MEM[22785];
assign MEM[29324] = MEM[22554] + MEM[22971];
assign MEM[29325] = MEM[22557] + MEM[22974];
assign MEM[29326] = MEM[22558] + MEM[22638];
assign MEM[29327] = MEM[22563] + MEM[22757];
assign MEM[29328] = MEM[22565] + MEM[22700];
assign MEM[29329] = MEM[22566] + MEM[22658];
assign MEM[29330] = MEM[22567] + MEM[22790];
assign MEM[29331] = MEM[22568] + MEM[22659];
assign MEM[29332] = MEM[22570] + MEM[22711];
assign MEM[29333] = MEM[22572] + MEM[22941];
assign MEM[29334] = MEM[22574] + MEM[22604];
assign MEM[29335] = MEM[22581] + MEM[24218];
assign MEM[29336] = MEM[22582] + MEM[22698];
assign MEM[29337] = MEM[22583] + MEM[22996];
assign MEM[29338] = MEM[22584] + MEM[22694];
assign MEM[29339] = MEM[22588] + MEM[22930];
assign MEM[29340] = MEM[22589] + MEM[23186];
assign MEM[29341] = MEM[22590] + MEM[22837];
assign MEM[29342] = MEM[22591] + MEM[23259];
assign MEM[29343] = MEM[22592] + MEM[23083];
assign MEM[29344] = MEM[22593] + MEM[22882];
assign MEM[29345] = MEM[22595] + MEM[22781];
assign MEM[29346] = MEM[22596] + MEM[22640];
assign MEM[29347] = MEM[22597] + MEM[22952];
assign MEM[29348] = MEM[22598] + MEM[23021];
assign MEM[29349] = MEM[22601] + MEM[24644];
assign MEM[29350] = MEM[22603] + MEM[22813];
assign MEM[29351] = MEM[22605] + MEM[24379];
assign MEM[29352] = MEM[22606] + MEM[22887];
assign MEM[29353] = MEM[22608] + MEM[22832];
assign MEM[29354] = MEM[22609] + MEM[22682];
assign MEM[29355] = MEM[22610] + MEM[23062];
assign MEM[29356] = MEM[22613] + MEM[22749];
assign MEM[29357] = MEM[22618] + MEM[22913];
assign MEM[29358] = MEM[22622] + MEM[22712];
assign MEM[29359] = MEM[22626] + MEM[23319];
assign MEM[29360] = MEM[22632] + MEM[22858];
assign MEM[29361] = MEM[22634] + MEM[22744];
assign MEM[29362] = MEM[22639] + MEM[22818];
assign MEM[29363] = MEM[22641] + MEM[22668];
assign MEM[29364] = MEM[22644] + MEM[22798];
assign MEM[29365] = MEM[22645] + MEM[22985];
assign MEM[29366] = MEM[22646] + MEM[23540];
assign MEM[29367] = MEM[22647] + MEM[24010];
assign MEM[29368] = MEM[22650] + MEM[22759];
assign MEM[29369] = MEM[22654] + MEM[23045];
assign MEM[29370] = MEM[22656] + MEM[22788];
assign MEM[29371] = MEM[22660] + MEM[23301];
assign MEM[29372] = MEM[22662] + MEM[22863];
assign MEM[29373] = MEM[22664] + MEM[22747];
assign MEM[29374] = MEM[22666] + MEM[22683];
assign MEM[29375] = MEM[22667] + MEM[22860];
assign MEM[29376] = MEM[22671] + MEM[22770];
assign MEM[29377] = MEM[22673] + MEM[22829];
assign MEM[29378] = MEM[22674] + MEM[23302];
assign MEM[29379] = MEM[22675] + MEM[22732];
assign MEM[29380] = MEM[22679] + MEM[22821];
assign MEM[29381] = MEM[22684] + MEM[22852];
assign MEM[29382] = MEM[22685] + MEM[22729];
assign MEM[29383] = MEM[22686] + MEM[22898];
assign MEM[29384] = MEM[22687] + MEM[22875];
assign MEM[29385] = MEM[22688] + MEM[22966];
assign MEM[29386] = MEM[22690] + MEM[22871];
assign MEM[29387] = MEM[22696] + MEM[22866];
assign MEM[29388] = MEM[22699] + MEM[23467];
assign MEM[29389] = MEM[22704] + MEM[22731];
assign MEM[29390] = MEM[22705] + MEM[22800];
assign MEM[29391] = MEM[22706] + MEM[22782];
assign MEM[29392] = MEM[22707] + MEM[22752];
assign MEM[29393] = MEM[22708] + MEM[22716];
assign MEM[29394] = MEM[22715] + MEM[22868];
assign MEM[29395] = MEM[22718] + MEM[23146];
assign MEM[29396] = MEM[22719] + MEM[24400];
assign MEM[29397] = MEM[22722] + MEM[22760];
assign MEM[29398] = MEM[22724] + MEM[23027];
assign MEM[29399] = MEM[22726] + MEM[22914];
assign MEM[29400] = MEM[22727] + MEM[22776];
assign MEM[29401] = MEM[22728] + MEM[23079];
assign MEM[29402] = MEM[22734] + MEM[23005];
assign MEM[29403] = MEM[22737] + MEM[22810];
assign MEM[29404] = MEM[22745] + MEM[23114];
assign MEM[29405] = MEM[22750] + MEM[22880];
assign MEM[29406] = MEM[22754] + MEM[23085];
assign MEM[29407] = MEM[22755] + MEM[22799];
assign MEM[29408] = MEM[22756] + MEM[22902];
assign MEM[29409] = MEM[22758] + MEM[23418];
assign MEM[29410] = MEM[22763] + MEM[22836];
assign MEM[29411] = MEM[22765] + MEM[23532];
assign MEM[29412] = MEM[22767] + MEM[22906];
assign MEM[29413] = MEM[22768] + MEM[23722];
assign MEM[29414] = MEM[22774] + MEM[23121];
assign MEM[29415] = MEM[22775] + MEM[22984];
assign MEM[29416] = MEM[22779] + MEM[23124];
assign MEM[29417] = MEM[22786] + MEM[23068];
assign MEM[29418] = MEM[22787] + MEM[23234];
assign MEM[29419] = MEM[22793] + MEM[23052];
assign MEM[29420] = MEM[22794] + MEM[22897];
assign MEM[29421] = MEM[22795] + MEM[23017];
assign MEM[29422] = MEM[22796] + MEM[22946];
assign MEM[29423] = MEM[22801] + MEM[23141];
assign MEM[29424] = MEM[22803] + MEM[23169];
assign MEM[29425] = MEM[22804] + MEM[23157];
assign MEM[29426] = MEM[22805] + MEM[23275];
assign MEM[29427] = MEM[22806] + MEM[23304];
assign MEM[29428] = MEM[22807] + MEM[23098];
assign MEM[29429] = MEM[22808] + MEM[23343];
assign MEM[29430] = MEM[22809] + MEM[24552];
assign MEM[29431] = MEM[22811] + MEM[22915];
assign MEM[29432] = MEM[22815] + MEM[24508];
assign MEM[29433] = MEM[22817] + MEM[22991];
assign MEM[29434] = MEM[22819] + MEM[22853];
assign MEM[29435] = MEM[22822] + MEM[23270];
assign MEM[29436] = MEM[22823] + MEM[22954];
assign MEM[29437] = MEM[22824] + MEM[23123];
assign MEM[29438] = MEM[22828] + MEM[23115];
assign MEM[29439] = MEM[22831] + MEM[22967];
assign MEM[29440] = MEM[22833] + MEM[22957];
assign MEM[29441] = MEM[22834] + MEM[23213];
assign MEM[29442] = MEM[22838] + MEM[23089];
assign MEM[29443] = MEM[22839] + MEM[23094];
assign MEM[29444] = MEM[22841] + MEM[23554];
assign MEM[29445] = MEM[22845] + MEM[23053];
assign MEM[29446] = MEM[22846] + MEM[22918];
assign MEM[29447] = MEM[22848] + MEM[23128];
assign MEM[29448] = MEM[22850] + MEM[22903];
assign MEM[29449] = MEM[22851] + MEM[22938];
assign MEM[29450] = MEM[22854] + MEM[23011];
assign MEM[29451] = MEM[22856] + MEM[22999];
assign MEM[29452] = MEM[22857] + MEM[23317];
assign MEM[29453] = MEM[22859] + MEM[23131];
assign MEM[29454] = MEM[22861] + MEM[22873];
assign MEM[29455] = MEM[22864] + MEM[23075];
assign MEM[29456] = MEM[22865] + MEM[23081];
assign MEM[29457] = MEM[22867] + MEM[23152];
assign MEM[29458] = MEM[22870] + MEM[22935];
assign MEM[29459] = MEM[22874] + MEM[23212];
assign MEM[29460] = MEM[22876] + MEM[22881];
assign MEM[29461] = MEM[22878] + MEM[23269];
assign MEM[29462] = MEM[22879] + MEM[24029];
assign MEM[29463] = MEM[22884] + MEM[23187];
assign MEM[29464] = MEM[22885] + MEM[23388];
assign MEM[29465] = MEM[22886] + MEM[22948];
assign MEM[29466] = MEM[22888] + MEM[24564];
assign MEM[29467] = MEM[22889] + MEM[23300];
assign MEM[29468] = MEM[22890] + MEM[22929];
assign MEM[29469] = MEM[22891] + MEM[23010];
assign MEM[29470] = MEM[22892] + MEM[23988];
assign MEM[29471] = MEM[22893] + MEM[23127];
assign MEM[29472] = MEM[22895] + MEM[23179];
assign MEM[29473] = MEM[22899] + MEM[23034];
assign MEM[29474] = MEM[22900] + MEM[23415];
assign MEM[29475] = MEM[22901] + MEM[23405];
assign MEM[29476] = MEM[22904] + MEM[23214];
assign MEM[29477] = MEM[22907] + MEM[23221];
assign MEM[29478] = MEM[22908] + MEM[23238];
assign MEM[29479] = MEM[22909] + MEM[23042];
assign MEM[29480] = MEM[22910] + MEM[24329];
assign MEM[29481] = MEM[22916] + MEM[23137];
assign MEM[29482] = MEM[22919] + MEM[23230];
assign MEM[29483] = MEM[22920] + MEM[23039];
assign MEM[29484] = MEM[22921] + MEM[22945];
assign MEM[29485] = MEM[22923] + MEM[23072];
assign MEM[29486] = MEM[22924] + MEM[24024];
assign MEM[29487] = MEM[22925] + MEM[23038];
assign MEM[29488] = MEM[22927] + MEM[22961];
assign MEM[29489] = MEM[22928] + MEM[22988];
assign MEM[29490] = MEM[22931] + MEM[23178];
assign MEM[29491] = MEM[22932] + MEM[23139];
assign MEM[29492] = MEM[22936] + MEM[23205];
assign MEM[29493] = MEM[22937] + MEM[22972];
assign MEM[29494] = MEM[22942] + MEM[22987];
assign MEM[29495] = MEM[22944] + MEM[23257];
assign MEM[29496] = MEM[22950] + MEM[23282];
assign MEM[29497] = MEM[22951] + MEM[23043];
assign MEM[29498] = MEM[22953] + MEM[23000];
assign MEM[29499] = MEM[22955] + MEM[23166];
assign MEM[29500] = MEM[22958] + MEM[23796];
assign MEM[29501] = MEM[22959] + MEM[23248];
assign MEM[29502] = MEM[22963] + MEM[23983];
assign MEM[29503] = MEM[22964] + MEM[23392];
assign MEM[29504] = MEM[22968] + MEM[23142];
assign MEM[29505] = MEM[22969] + MEM[23480];
assign MEM[29506] = MEM[22970] + MEM[23057];
assign MEM[29507] = MEM[22973] + MEM[24943];
assign MEM[29508] = MEM[22975] + MEM[24208];
assign MEM[29509] = MEM[22976] + MEM[23070];
assign MEM[29510] = MEM[22977] + MEM[23035];
assign MEM[29511] = MEM[22978] + MEM[23315];
assign MEM[29512] = MEM[22980] + MEM[23134];
assign MEM[29513] = MEM[22981] + MEM[23742];
assign MEM[29514] = MEM[22982] + MEM[23076];
assign MEM[29515] = MEM[22983] + MEM[23140];
assign MEM[29516] = MEM[22986] + MEM[23087];
assign MEM[29517] = MEM[22989] + MEM[23080];
assign MEM[29518] = MEM[22990] + MEM[23051];
assign MEM[29519] = MEM[22992] + MEM[23231];
assign MEM[29520] = MEM[22993] + MEM[23008];
assign MEM[29521] = MEM[22994] + MEM[23426];
assign MEM[29522] = MEM[22995] + MEM[23761];
assign MEM[29523] = MEM[22997] + MEM[23245];
assign MEM[29524] = MEM[22998] + MEM[23402];
assign MEM[29525] = MEM[23001] + MEM[23028];
assign MEM[29526] = MEM[23002] + MEM[23096];
assign MEM[29527] = MEM[23003] + MEM[23328];
assign MEM[29528] = MEM[23004] + MEM[23326];
assign MEM[29529] = MEM[23006] + MEM[23965];
assign MEM[29530] = MEM[23009] + MEM[23036];
assign MEM[29531] = MEM[23012] + MEM[23784];
assign MEM[29532] = MEM[23013] + MEM[23119];
assign MEM[29533] = MEM[23014] + MEM[23180];
assign MEM[29534] = MEM[23015] + MEM[23258];
assign MEM[29535] = MEM[23016] + MEM[23250];
assign MEM[29536] = MEM[23019] + MEM[23336];
assign MEM[29537] = MEM[23024] + MEM[23279];
assign MEM[29538] = MEM[23026] + MEM[23543];
assign MEM[29539] = MEM[23029] + MEM[23144];
assign MEM[29540] = MEM[23031] + MEM[23577];
assign MEM[29541] = MEM[23032] + MEM[23159];
assign MEM[29542] = MEM[23033] + MEM[23165];
assign MEM[29543] = MEM[23037] + MEM[23277];
assign MEM[29544] = MEM[23040] + MEM[23756];
assign MEM[29545] = MEM[23041] + MEM[23046];
assign MEM[29546] = MEM[23044] + MEM[23067];
assign MEM[29547] = MEM[23048] + MEM[23078];
assign MEM[29548] = MEM[23049] + MEM[23284];
assign MEM[29549] = MEM[23050] + MEM[24433];
assign MEM[29550] = MEM[23054] + MEM[23314];
assign MEM[29551] = MEM[23055] + MEM[23104];
assign MEM[29552] = MEM[23056] + MEM[23265];
assign MEM[29553] = MEM[23058] + MEM[23737];
assign MEM[29554] = MEM[23060] + MEM[23160];
assign MEM[29555] = MEM[23061] + MEM[23646];
assign MEM[29556] = MEM[23063] + MEM[23609];
assign MEM[29557] = MEM[23064] + MEM[23066];
assign MEM[29558] = MEM[23065] + MEM[23111];
assign MEM[29559] = MEM[23069] + MEM[23979];
assign MEM[29560] = MEM[23071] + MEM[23185];
assign MEM[29561] = MEM[23073] + MEM[23138];
assign MEM[29562] = MEM[23074] + MEM[23501];
assign MEM[29563] = MEM[23077] + MEM[23154];
assign MEM[29564] = MEM[23082] + MEM[23202];
assign MEM[29565] = MEM[23084] + MEM[23586];
assign MEM[29566] = MEM[23086] + MEM[24958];
assign MEM[29567] = MEM[23088] + MEM[23091];
assign MEM[29568] = MEM[23092] + MEM[23135];
assign MEM[29569] = MEM[23093] + MEM[23246];
assign MEM[29570] = MEM[23095] + MEM[23145];
assign MEM[29571] = MEM[23097] + MEM[23690];
assign MEM[29572] = MEM[23099] + MEM[23892];
assign MEM[29573] = MEM[23100] + MEM[23174];
assign MEM[29574] = MEM[23101] + MEM[24510];
assign MEM[29575] = MEM[23102] + MEM[23359];
assign MEM[29576] = MEM[23103] + MEM[23266];
assign MEM[29577] = MEM[23106] + MEM[24451];
assign MEM[29578] = MEM[23107] + MEM[23339];
assign MEM[29579] = MEM[23108] + MEM[23183];
assign MEM[29580] = MEM[23109] + MEM[23227];
assign MEM[29581] = MEM[23110] + MEM[23893];
assign MEM[29582] = MEM[23112] + MEM[23453];
assign MEM[29583] = MEM[23113] + MEM[24469];
assign MEM[29584] = MEM[23116] + MEM[23161];
assign MEM[29585] = MEM[23120] + MEM[23182];
assign MEM[29586] = MEM[23125] + MEM[23253];
assign MEM[29587] = MEM[23126] + MEM[24677];
assign MEM[29588] = MEM[23130] + MEM[23313];
assign MEM[29589] = MEM[23132] + MEM[24733];
assign MEM[29590] = MEM[23133] + MEM[23341];
assign MEM[29591] = MEM[23136] + MEM[23271];
assign MEM[29592] = MEM[23143] + MEM[23170];
assign MEM[29593] = MEM[23147] + MEM[23872];
assign MEM[29594] = MEM[23148] + MEM[23377];
assign MEM[29595] = MEM[23149] + MEM[24097];
assign MEM[29596] = MEM[23150] + MEM[23307];
assign MEM[29597] = MEM[23151] + MEM[24425];
assign MEM[29598] = MEM[23153] + MEM[23946];
assign MEM[29599] = MEM[23156] + MEM[23472];
assign MEM[29600] = MEM[23158] + MEM[24277];
assign MEM[29601] = MEM[23163] + MEM[23176];
assign MEM[29602] = MEM[23164] + MEM[23200];
assign MEM[29603] = MEM[23167] + MEM[24173];
assign MEM[29604] = MEM[23168] + MEM[23236];
assign MEM[29605] = MEM[23171] + MEM[23475];
assign MEM[29606] = MEM[23172] + MEM[23972];
assign MEM[29607] = MEM[23173] + MEM[23192];
assign MEM[29608] = MEM[23175] + MEM[23184];
assign MEM[29609] = MEM[23177] + MEM[23324];
assign MEM[29610] = MEM[23181] + MEM[23303];
assign MEM[29611] = MEM[23188] + MEM[23261];
assign MEM[29612] = MEM[23189] + MEM[23631];
assign MEM[29613] = MEM[23190] + MEM[23241];
assign MEM[29614] = MEM[23191] + MEM[23349];
assign MEM[29615] = MEM[23193] + MEM[23397];
assign MEM[29616] = MEM[23194] + MEM[23375];
assign MEM[29617] = MEM[23195] + MEM[23207];
assign MEM[29618] = MEM[23196] + MEM[23360];
assign MEM[29619] = MEM[23198] + MEM[24153];
assign MEM[29620] = MEM[23199] + MEM[24078];
assign MEM[29621] = MEM[23201] + MEM[23505];
assign MEM[29622] = MEM[23203] + MEM[23461];
assign MEM[29623] = MEM[23204] + MEM[24566];
assign MEM[29624] = MEM[23206] + MEM[24654];
assign MEM[29625] = MEM[23208] + MEM[23263];
assign MEM[29626] = MEM[23209] + MEM[23476];
assign MEM[29627] = MEM[23210] + MEM[23229];
assign MEM[29628] = MEM[23211] + MEM[23260];
assign MEM[29629] = MEM[23215] + MEM[23254];
assign MEM[29630] = MEM[23216] + MEM[23267];
assign MEM[29631] = MEM[23217] + MEM[23308];
assign MEM[29632] = MEM[23218] + MEM[23237];
assign MEM[29633] = MEM[23219] + MEM[23803];
assign MEM[29634] = MEM[23220] + MEM[23247];
assign MEM[29635] = MEM[23222] + MEM[23985];
assign MEM[29636] = MEM[23223] + MEM[23327];
assign MEM[29637] = MEM[23224] + MEM[23922];
assign MEM[29638] = MEM[23225] + MEM[23529];
assign MEM[29639] = MEM[23226] + MEM[23450];
assign MEM[29640] = MEM[23228] + MEM[23340];
assign MEM[29641] = MEM[23232] + MEM[23443];
assign MEM[29642] = MEM[23233] + MEM[24357];
assign MEM[29643] = MEM[23235] + MEM[23290];
assign MEM[29644] = MEM[23239] + MEM[23466];
assign MEM[29645] = MEM[23240] + MEM[23484];
assign MEM[29646] = MEM[23242] + MEM[23527];
assign MEM[29647] = MEM[23244] + MEM[23305];
assign MEM[29648] = MEM[23249] + MEM[24125];
assign MEM[29649] = MEM[23251] + MEM[23499];
assign MEM[29650] = MEM[23252] + MEM[23481];
assign MEM[29651] = MEM[23255] + MEM[23731];
assign MEM[29652] = MEM[23256] + MEM[23346];
assign MEM[29653] = MEM[23262] + MEM[23347];
assign MEM[29654] = MEM[23264] + MEM[24611];
assign MEM[29655] = MEM[23268] + MEM[23664];
assign MEM[29656] = MEM[23272] + MEM[23750];
assign MEM[29657] = MEM[23273] + MEM[24612];
assign MEM[29658] = MEM[23276] + MEM[24307];
assign MEM[29659] = MEM[23278] + MEM[23486];
assign MEM[29660] = MEM[23280] + MEM[23350];
assign MEM[29661] = MEM[23281] + MEM[23353];
assign MEM[29662] = MEM[23283] + MEM[23358];
assign MEM[29663] = MEM[23285] + MEM[23356];
assign MEM[29664] = MEM[23286] + MEM[24107];
assign MEM[29665] = MEM[23287] + MEM[23296];
assign MEM[29666] = MEM[23288] + MEM[23292];
assign MEM[29667] = MEM[23289] + MEM[23624];
assign MEM[29668] = MEM[23291] + MEM[24298];
assign MEM[29669] = MEM[23293] + MEM[24018];
assign MEM[29670] = MEM[23294] + MEM[24025];
assign MEM[29671] = MEM[23295] + MEM[23535];
assign MEM[29672] = MEM[23297] + MEM[23478];
assign MEM[29673] = MEM[23298] + MEM[24891];
assign MEM[29674] = MEM[23299] + MEM[23396];
assign MEM[29675] = MEM[23306] + MEM[23864];
assign MEM[29676] = MEM[23309] + MEM[23982];
assign MEM[29677] = MEM[23311] + MEM[23623];
assign MEM[29678] = MEM[23312] + MEM[24286];
assign MEM[29679] = MEM[23316] + MEM[24028];
assign MEM[29680] = MEM[23318] + MEM[23545];
assign MEM[29681] = MEM[23320] + MEM[23458];
assign MEM[29682] = MEM[23321] + MEM[23510];
assign MEM[29683] = MEM[23322] + MEM[24004];
assign MEM[29684] = MEM[23323] + MEM[23560];
assign MEM[29685] = MEM[23325] + MEM[23464];
assign MEM[29686] = MEM[23329] + MEM[23878];
assign MEM[29687] = MEM[23330] + MEM[23820];
assign MEM[29688] = MEM[23331] + MEM[24637];
assign MEM[29689] = MEM[23332] + MEM[23628];
assign MEM[29690] = MEM[23333] + MEM[23615];
assign MEM[29691] = MEM[23334] + MEM[24386];
assign MEM[29692] = MEM[23335] + MEM[24086];
assign MEM[29693] = MEM[23337] + MEM[23593];
assign MEM[29694] = MEM[23338] + MEM[23821];
assign MEM[29695] = MEM[23342] + MEM[24013];
assign MEM[29696] = MEM[23344] + MEM[24043];
assign MEM[29697] = MEM[23345] + MEM[24559];
assign MEM[29698] = MEM[23351] + MEM[23367];
assign MEM[29699] = MEM[23352] + MEM[24030];
assign MEM[29700] = MEM[23354] + MEM[24498];
assign MEM[29701] = MEM[23355] + MEM[23368];
assign MEM[29702] = MEM[23357] + MEM[23611];
assign MEM[29703] = MEM[23361] + MEM[24624];
assign MEM[29704] = MEM[23362] + MEM[23826];
assign MEM[29705] = MEM[23363] + MEM[24299];
assign MEM[29706] = MEM[23364] + MEM[23942];
assign MEM[29707] = MEM[23365] + MEM[25126];
assign MEM[29708] = MEM[23369] + MEM[27060];
assign MEM[29709] = MEM[23370] + MEM[26478];
assign MEM[29710] = MEM[23371] + MEM[24944];
assign MEM[29711] = MEM[23372] + MEM[24853];
assign MEM[29712] = MEM[23373] + MEM[24631];
assign MEM[29713] = MEM[23374] + MEM[26769];
assign MEM[29714] = MEM[23376] + MEM[24439];
assign MEM[29715] = MEM[23378] + MEM[24068];
assign MEM[29716] = MEM[23379] + MEM[24860];
assign MEM[29717] = MEM[23380] + MEM[24623];
assign MEM[29718] = MEM[23381] + MEM[24441];
assign MEM[29719] = MEM[23382] + MEM[25757];
assign MEM[29720] = MEM[23383] + MEM[25402];
assign MEM[29721] = MEM[23384] + MEM[24591];
assign MEM[29722] = MEM[23385] + MEM[29308];
assign MEM[29723] = MEM[23386] + MEM[25817];
assign MEM[29724] = MEM[23387] + MEM[28443];
assign MEM[29725] = MEM[23389] + MEM[24966];
assign MEM[29726] = MEM[23390] + MEM[26459];
assign MEM[29727] = MEM[23393] + MEM[25911];
assign MEM[29728] = MEM[23394] + MEM[26127];
assign MEM[29729] = MEM[23395] + MEM[23825];
assign MEM[29730] = MEM[23398] + MEM[26099];
assign MEM[29731] = MEM[23399] + MEM[24832];
assign MEM[29732] = MEM[23400] + MEM[24918];
assign MEM[29733] = MEM[23401] + MEM[29236];
assign MEM[29734] = MEM[23403] + MEM[23641];
assign MEM[29735] = MEM[23404] + MEM[26836];
assign MEM[29736] = MEM[23406] + MEM[23728];
assign MEM[29737] = MEM[23407] + MEM[28102];
assign MEM[29738] = MEM[23408] + MEM[24283];
assign MEM[29739] = MEM[23409] + MEM[24968];
assign MEM[29740] = MEM[23410] + MEM[24333];
assign MEM[29741] = MEM[23411] + MEM[24594];
assign MEM[29742] = MEM[23412] + MEM[25362];
assign MEM[29743] = MEM[23413] + MEM[24487];
assign MEM[29744] = MEM[23414] + MEM[25474];
assign MEM[29745] = MEM[23416] + MEM[26081];
assign MEM[29746] = MEM[23417] + MEM[26978];
assign MEM[29747] = MEM[23419] + MEM[26029];
assign MEM[29748] = MEM[23420] + MEM[24738];
assign MEM[29749] = MEM[23421] + MEM[25452];
assign MEM[29750] = MEM[23422] + MEM[26274];
assign MEM[29751] = MEM[23423] + MEM[23512];
assign MEM[29752] = MEM[23424] + MEM[24807];
assign MEM[29753] = MEM[23425] + MEM[23963];
assign MEM[29754] = MEM[23427] + MEM[24335];
assign MEM[29755] = MEM[23428] + MEM[23619];
assign MEM[29756] = MEM[23429] + MEM[23842];
assign MEM[29757] = MEM[23431] + MEM[25198];
assign MEM[29758] = MEM[23432] + MEM[24534];
assign MEM[29759] = MEM[23433] + MEM[24695];
assign MEM[29760] = MEM[23434] + MEM[23700];
assign MEM[29761] = MEM[23435] + MEM[25284];
assign MEM[29762] = MEM[23436] + MEM[24609];
assign MEM[29763] = MEM[23437] + MEM[25186];
assign MEM[29764] = MEM[23438] + MEM[25352];
assign MEM[29765] = MEM[23439] + MEM[28809];
assign MEM[29766] = MEM[23440] + MEM[24574];
assign MEM[29767] = MEM[23441] + MEM[23871];
assign MEM[29768] = MEM[23442] + MEM[27737];
assign MEM[29769] = MEM[23444] + MEM[25470];
assign MEM[29770] = MEM[23445] + MEM[26406];
assign MEM[29771] = MEM[23446] + MEM[25334];
assign MEM[29772] = MEM[23447] + MEM[24124];
assign MEM[29773] = MEM[23448] + MEM[26526];
assign MEM[29774] = MEM[23449] + MEM[25336];
assign MEM[29775] = MEM[23451] + MEM[25009];
assign MEM[29776] = MEM[23452] + MEM[26119];
assign MEM[29777] = MEM[23454] + MEM[25209];
assign MEM[29778] = MEM[23455] + MEM[28529];
assign MEM[29779] = MEM[23456] + MEM[25865];
assign MEM[29780] = MEM[23459] + MEM[25428];
assign MEM[29781] = MEM[23460] + MEM[25028];
assign MEM[29782] = MEM[23462] + MEM[29142];
assign MEM[29783] = MEM[23463] + MEM[23808];
assign MEM[29784] = MEM[23465] + MEM[25732];
assign MEM[29785] = MEM[23468] + MEM[24717];
assign MEM[29786] = MEM[23469] + MEM[27016];
assign MEM[29787] = MEM[23470] + MEM[24914];
assign MEM[29788] = MEM[23471] + MEM[29362];
assign MEM[29789] = MEM[23473] + MEM[25810];
assign MEM[29790] = MEM[23474] + MEM[25589];
assign MEM[29791] = MEM[23477] + MEM[25856];
assign MEM[29792] = MEM[23479] + MEM[24026];
assign MEM[29793] = MEM[23482] + MEM[28164];
assign MEM[29794] = MEM[23483] + MEM[25801];
assign MEM[29795] = MEM[23485] + MEM[26999];
assign MEM[29796] = MEM[23488] + MEM[24461];
assign MEM[29797] = MEM[23489] + MEM[27979];
assign MEM[29798] = MEM[23490] + MEM[25374];
assign MEM[29799] = MEM[23491] + MEM[26143];
assign MEM[29800] = MEM[23492] + MEM[25747];
assign MEM[29801] = MEM[23493] + MEM[26087];
assign MEM[29802] = MEM[23494] + MEM[25588];
assign MEM[29803] = MEM[23495] + MEM[26370];
assign MEM[29804] = MEM[23496] + MEM[24099];
assign MEM[29805] = MEM[23497] + MEM[26874];
assign MEM[29806] = MEM[23498] + MEM[27320];
assign MEM[29807] = MEM[23500] + MEM[25003];
assign MEM[29808] = MEM[23502] + MEM[23754];
assign MEM[29809] = MEM[23503] + MEM[24587];
assign MEM[29810] = MEM[23504] + MEM[24529];
assign MEM[29811] = MEM[23506] + MEM[29329];
assign MEM[29812] = MEM[23507] + MEM[26808];
assign MEM[29813] = MEM[23508] + MEM[24744];
assign MEM[29814] = MEM[23509] + MEM[29372];
assign MEM[29815] = MEM[23511] + MEM[24814];
assign MEM[29816] = MEM[23513] + MEM[24697];
assign MEM[29817] = MEM[23514] + MEM[25121];
assign MEM[29818] = MEM[23515] + MEM[25597];
assign MEM[29819] = MEM[23516] + MEM[24685];
assign MEM[29820] = MEM[23517] + MEM[24232];
assign MEM[29821] = MEM[23518] + MEM[25957];
assign MEM[29822] = MEM[23519] + MEM[25825];
assign MEM[29823] = MEM[23520] + MEM[25033];
assign MEM[29824] = MEM[23521] + MEM[26170];
assign MEM[29825] = MEM[23522] + MEM[25699];
assign MEM[29826] = MEM[23523] + MEM[24823];
assign MEM[29827] = MEM[23524] + MEM[24785];
assign MEM[29828] = MEM[23525] + MEM[24505];
assign MEM[29829] = MEM[23526] + MEM[27193];
assign MEM[29830] = MEM[23528] + MEM[26831];
assign MEM[29831] = MEM[23531] + MEM[23907];
assign MEM[29832] = MEM[23533] + MEM[25380];
assign MEM[29833] = MEM[23534] + MEM[26785];
assign MEM[29834] = MEM[23536] + MEM[25901];
assign MEM[29835] = MEM[23537] + MEM[23695];
assign MEM[29836] = MEM[23538] + MEM[23726];
assign MEM[29837] = MEM[23539] + MEM[24845];
assign MEM[29838] = MEM[23541] + MEM[24061];
assign MEM[29839] = MEM[23542] + MEM[26488];
assign MEM[29840] = MEM[23544] + MEM[25715];
assign MEM[29841] = MEM[23546] + MEM[25656];
assign MEM[29842] = MEM[23547] + MEM[25999];
assign MEM[29843] = MEM[23548] + MEM[23758];
assign MEM[29844] = MEM[23549] + MEM[25375];
assign MEM[29845] = MEM[23550] + MEM[24841];
assign MEM[29846] = MEM[23551] + MEM[25413];
assign MEM[29847] = MEM[23552] + MEM[29031];
assign MEM[29848] = MEM[23553] + MEM[26545];
assign MEM[29849] = MEM[23555] + MEM[25298];
assign MEM[29850] = MEM[23556] + MEM[25176];
assign MEM[29851] = MEM[23557] + MEM[24409];
assign MEM[29852] = MEM[23559] + MEM[25257];
assign MEM[29853] = MEM[23561] + MEM[24652];
assign MEM[29854] = MEM[23562] + MEM[24122];
assign MEM[29855] = MEM[23563] + MEM[25165];
assign MEM[29856] = MEM[23564] + MEM[24150];
assign MEM[29857] = MEM[23565] + MEM[27214];
assign MEM[29858] = MEM[23566] + MEM[24893];
assign MEM[29859] = MEM[23567] + MEM[24514];
assign MEM[29860] = MEM[23568] + MEM[24758];
assign MEM[29861] = MEM[23569] + MEM[24795];
assign MEM[29862] = MEM[23570] + MEM[24364];
assign MEM[29863] = MEM[23571] + MEM[26438];
assign MEM[29864] = MEM[23572] + MEM[25169];
assign MEM[29865] = MEM[23573] + MEM[24867];
assign MEM[29866] = MEM[23574] + MEM[24511];
assign MEM[29867] = MEM[23575] + MEM[24694];
assign MEM[29868] = MEM[23576] + MEM[24290];
assign MEM[29869] = MEM[23578] + MEM[26610];
assign MEM[29870] = MEM[23579] + MEM[27218];
assign MEM[29871] = MEM[23580] + MEM[24641];
assign MEM[29872] = MEM[23581] + MEM[24635];
assign MEM[29873] = MEM[23582] + MEM[27126];
assign MEM[29874] = MEM[23583] + MEM[26223];
assign MEM[29875] = MEM[23584] + MEM[24597];
assign MEM[29876] = MEM[23585] + MEM[26516];
assign MEM[29877] = MEM[23587] + MEM[27034];
assign MEM[29878] = MEM[23588] + MEM[28626];
assign MEM[29879] = MEM[23589] + MEM[25695];
assign MEM[29880] = MEM[23590] + MEM[25061];
assign MEM[29881] = MEM[23591] + MEM[25490];
assign MEM[29882] = MEM[23592] + MEM[25816];
assign MEM[29883] = MEM[23594] + MEM[24447];
assign MEM[29884] = MEM[23595] + MEM[24321];
assign MEM[29885] = MEM[23596] + MEM[28049];
assign MEM[29886] = MEM[23597] + MEM[28422];
assign MEM[29887] = MEM[23598] + MEM[25861];
assign MEM[29888] = MEM[23599] + MEM[27572];
assign MEM[29889] = MEM[23600] + MEM[27516];
assign MEM[29890] = MEM[23601] + MEM[25060];
assign MEM[29891] = MEM[23602] + MEM[27261];
assign MEM[29892] = MEM[23603] + MEM[24359];
assign MEM[29893] = MEM[23604] + MEM[24957];
assign MEM[29894] = MEM[23605] + MEM[25201];
assign MEM[29895] = MEM[23606] + MEM[25776];
assign MEM[29896] = MEM[23607] + MEM[25814];
assign MEM[29897] = MEM[23608] + MEM[27339];
assign MEM[29898] = MEM[23610] + MEM[24166];
assign MEM[29899] = MEM[23612] + MEM[24523];
assign MEM[29900] = MEM[23613] + MEM[24788];
assign MEM[29901] = MEM[23614] + MEM[23924];
assign MEM[29902] = MEM[23616] + MEM[26012];
assign MEM[29903] = MEM[23617] + MEM[25150];
assign MEM[29904] = MEM[23618] + MEM[27078];
assign MEM[29905] = MEM[23620] + MEM[25722];
assign MEM[29906] = MEM[23621] + MEM[25379];
assign MEM[29907] = MEM[23622] + MEM[26704];
assign MEM[29908] = MEM[23625] + MEM[26604];
assign MEM[29909] = MEM[23626] + MEM[25238];
assign MEM[29910] = MEM[23627] + MEM[23823];
assign MEM[29911] = MEM[23629] + MEM[26091];
assign MEM[29912] = MEM[23630] + MEM[25812];
assign MEM[29913] = MEM[23632] + MEM[25012];
assign MEM[29914] = MEM[23633] + MEM[26702];
assign MEM[29915] = MEM[23634] + MEM[24032];
assign MEM[29916] = MEM[23635] + MEM[26366];
assign MEM[29917] = MEM[23636] + MEM[24203];
assign MEM[29918] = MEM[23637] + MEM[24797];
assign MEM[29919] = MEM[23638] + MEM[25044];
assign MEM[29920] = MEM[23639] + MEM[26612];
assign MEM[29921] = MEM[23640] + MEM[25743];
assign MEM[29922] = MEM[23642] + MEM[24223];
assign MEM[29923] = MEM[23643] + MEM[27127];
assign MEM[29924] = MEM[23644] + MEM[26758];
assign MEM[29925] = MEM[23645] + MEM[25275];
assign MEM[29926] = MEM[23647] + MEM[24391];
assign MEM[29927] = MEM[23648] + MEM[25129];
assign MEM[29928] = MEM[23649] + MEM[23930];
assign MEM[29929] = MEM[23650] + MEM[25382];
assign MEM[29930] = MEM[23651] + MEM[27304];
assign MEM[29931] = MEM[23652] + MEM[27148];
assign MEM[29932] = MEM[23653] + MEM[26324];
assign MEM[29933] = MEM[23654] + MEM[28523];
assign MEM[29934] = MEM[23655] + MEM[24296];
assign MEM[29935] = MEM[23656] + MEM[26980];
assign MEM[29936] = MEM[23657] + MEM[25187];
assign MEM[29937] = MEM[23658] + MEM[24761];
assign MEM[29938] = MEM[23660] + MEM[27322];
assign MEM[29939] = MEM[23661] + MEM[25270];
assign MEM[29940] = MEM[23662] + MEM[28972];
assign MEM[29941] = MEM[23663] + MEM[25195];
assign MEM[29942] = MEM[23665] + MEM[25410];
assign MEM[29943] = MEM[23666] + MEM[25500];
assign MEM[29944] = MEM[23667] + MEM[25024];
assign MEM[29945] = MEM[23668] + MEM[24317];
assign MEM[29946] = MEM[23669] + MEM[24656];
assign MEM[29947] = MEM[23670] + MEM[25727];
assign MEM[29948] = MEM[23671] + MEM[25744];
assign MEM[29949] = MEM[23672] + MEM[25389];
assign MEM[29950] = MEM[23673] + MEM[25055];
assign MEM[29951] = MEM[23674] + MEM[27093];
assign MEM[29952] = MEM[23675] + MEM[24116];
assign MEM[29953] = MEM[23676] + MEM[25149];
assign MEM[29954] = MEM[23677] + MEM[24667];
assign MEM[29955] = MEM[23678] + MEM[24464];
assign MEM[29956] = MEM[23679] + MEM[28019];
assign MEM[29957] = MEM[23680] + MEM[24521];
assign MEM[29958] = MEM[23681] + MEM[26484];
assign MEM[29959] = MEM[23682] + MEM[24438];
assign MEM[29960] = MEM[23683] + MEM[25842];
assign MEM[29961] = MEM[23686] + MEM[24353];
assign MEM[29962] = MEM[23687] + MEM[26664];
assign MEM[29963] = MEM[23688] + MEM[26354];
assign MEM[29964] = MEM[23689] + MEM[25035];
assign MEM[29965] = MEM[23691] + MEM[26130];
assign MEM[29966] = MEM[23692] + MEM[24872];
assign MEM[29967] = MEM[23693] + MEM[25276];
assign MEM[29968] = MEM[23694] + MEM[25163];
assign MEM[29969] = MEM[23696] + MEM[25366];
assign MEM[29970] = MEM[23697] + MEM[27902];
assign MEM[29971] = MEM[23698] + MEM[25910];
assign MEM[29972] = MEM[23699] + MEM[24782];
assign MEM[29973] = MEM[23701] + MEM[24712];
assign MEM[29974] = MEM[23702] + MEM[25089];
assign MEM[29975] = MEM[23703] + MEM[24729];
assign MEM[29976] = MEM[23704] + MEM[25233];
assign MEM[29977] = MEM[23705] + MEM[24370];
assign MEM[29978] = MEM[23706] + MEM[26590];
assign MEM[29979] = MEM[23707] + MEM[29346];
assign MEM[29980] = MEM[23708] + MEM[25037];
assign MEM[29981] = MEM[23709] + MEM[24497];
assign MEM[29982] = MEM[23710] + MEM[27992];
assign MEM[29983] = MEM[23711] + MEM[25192];
assign MEM[29984] = MEM[23712] + MEM[25502];
assign MEM[29985] = MEM[23713] + MEM[26804];
assign MEM[29986] = MEM[23714] + MEM[28160];
assign MEM[29987] = MEM[23716] + MEM[24202];
assign MEM[29988] = MEM[23717] + MEM[24555];
assign MEM[29989] = MEM[23718] + MEM[24750];
assign MEM[29990] = MEM[23719] + MEM[28985];
assign MEM[29991] = MEM[23720] + MEM[29645];
assign MEM[29992] = MEM[23721] + MEM[23863];
assign MEM[29993] = MEM[23723] + MEM[28642];
assign MEM[29994] = MEM[23724] + MEM[25730];
assign MEM[29995] = MEM[23725] + MEM[26499];
assign MEM[29996] = MEM[23727] + MEM[24897];
assign MEM[29997] = MEM[23729] + MEM[24426];
assign MEM[29998] = MEM[23730] + MEM[26110];
assign MEM[29999] = MEM[23732] + MEM[25119];
assign MEM[30000] = MEM[23733] + MEM[25506];
assign MEM[30001] = MEM[23734] + MEM[25311];
assign MEM[30002] = MEM[23735] + MEM[24027];
assign MEM[30003] = MEM[23736] + MEM[24820];
assign MEM[30004] = MEM[23738] + MEM[25606];
assign MEM[30005] = MEM[23739] + MEM[25648];
assign MEM[30006] = MEM[23740] + MEM[24374];
assign MEM[30007] = MEM[23741] + MEM[24481];
assign MEM[30008] = MEM[23743] + MEM[24870];
assign MEM[30009] = MEM[23744] + MEM[25923];
assign MEM[30010] = MEM[23745] + MEM[25881];
assign MEM[30011] = MEM[23746] + MEM[24809];
assign MEM[30012] = MEM[23747] + MEM[24843];
assign MEM[30013] = MEM[23748] + MEM[25248];
assign MEM[30014] = MEM[23749] + MEM[24741];
assign MEM[30015] = MEM[23751] + MEM[23769];
assign MEM[30016] = MEM[23752] + MEM[24181];
assign MEM[30017] = MEM[23753] + MEM[25745];
assign MEM[30018] = MEM[23755] + MEM[24349];
assign MEM[30019] = MEM[23757] + MEM[26123];
assign MEM[30020] = MEM[23760] + MEM[24948];
assign MEM[30021] = MEM[23763] + MEM[24198];
assign MEM[30022] = MEM[23764] + MEM[28444];
assign MEM[30023] = MEM[23765] + MEM[24996];
assign MEM[30024] = MEM[23766] + MEM[24524];
assign MEM[30025] = MEM[23767] + MEM[25967];
assign MEM[30026] = MEM[23768] + MEM[25593];
assign MEM[30027] = MEM[23770] + MEM[26689];
assign MEM[30028] = MEM[23771] + MEM[24680];
assign MEM[30029] = MEM[23772] + MEM[28087];
assign MEM[30030] = MEM[23773] + MEM[24162];
assign MEM[30031] = MEM[23774] + MEM[24813];
assign MEM[30032] = MEM[23775] + MEM[25053];
assign MEM[30033] = MEM[23776] + MEM[25364];
assign MEM[30034] = MEM[23777] + MEM[25016];
assign MEM[30035] = MEM[23778] + MEM[25054];
assign MEM[30036] = MEM[23779] + MEM[25237];
assign MEM[30037] = MEM[23780] + MEM[24900];
assign MEM[30038] = MEM[23781] + MEM[24619];
assign MEM[30039] = MEM[23782] + MEM[24268];
assign MEM[30040] = MEM[23783] + MEM[24976];
assign MEM[30041] = MEM[23785] + MEM[26013];
assign MEM[30042] = MEM[23786] + MEM[24734];
assign MEM[30043] = MEM[23787] + MEM[24790];
assign MEM[30044] = MEM[23788] + MEM[25207];
assign MEM[30045] = MEM[23789] + MEM[25558];
assign MEM[30046] = MEM[23790] + MEM[26311];
assign MEM[30047] = MEM[23791] + MEM[27788];
assign MEM[30048] = MEM[23792] + MEM[26383];
assign MEM[30049] = MEM[23793] + MEM[28442];
assign MEM[30050] = MEM[23794] + MEM[24052];
assign MEM[30051] = MEM[23795] + MEM[26073];
assign MEM[30052] = MEM[23797] + MEM[25676];
assign MEM[30053] = MEM[23798] + MEM[24940];
assign MEM[30054] = MEM[23799] + MEM[25711];
assign MEM[30055] = MEM[23800] + MEM[25032];
assign MEM[30056] = MEM[23801] + MEM[26555];
assign MEM[30057] = MEM[23802] + MEM[24852];
assign MEM[30058] = MEM[23804] + MEM[24323];
assign MEM[30059] = MEM[23806] + MEM[24647];
assign MEM[30060] = MEM[23807] + MEM[25437];
assign MEM[30061] = MEM[23809] + MEM[27298];
assign MEM[30062] = MEM[23810] + MEM[24875];
assign MEM[30063] = MEM[23811] + MEM[26443];
assign MEM[30064] = MEM[23812] + MEM[24460];
assign MEM[30065] = MEM[23813] + MEM[24221];
assign MEM[30066] = MEM[23814] + MEM[25418];
assign MEM[30067] = MEM[23815] + MEM[28715];
assign MEM[30068] = MEM[23816] + MEM[24678];
assign MEM[30069] = MEM[23817] + MEM[26175];
assign MEM[30070] = MEM[23818] + MEM[25976];
assign MEM[30071] = MEM[23819] + MEM[24686];
assign MEM[30072] = MEM[23822] + MEM[24925];
assign MEM[30073] = MEM[23824] + MEM[26009];
assign MEM[30074] = MEM[23827] + MEM[27069];
assign MEM[30075] = MEM[23828] + MEM[28865];
assign MEM[30076] = MEM[23830] + MEM[24551];
assign MEM[30077] = MEM[23831] + MEM[24408];
assign MEM[30078] = MEM[23832] + MEM[26811];
assign MEM[30079] = MEM[23833] + MEM[26525];
assign MEM[30080] = MEM[23834] + MEM[25125];
assign MEM[30081] = MEM[23835] + MEM[24186];
assign MEM[30082] = MEM[23836] + MEM[25719];
assign MEM[30083] = MEM[23837] + MEM[26523];
assign MEM[30084] = MEM[23838] + MEM[23841];
assign MEM[30085] = MEM[23839] + MEM[25914];
assign MEM[30086] = MEM[23840] + MEM[24868];
assign MEM[30087] = MEM[23843] + MEM[24557];
assign MEM[30088] = MEM[23844] + MEM[26113];
assign MEM[30089] = MEM[23845] + MEM[27019];
assign MEM[30090] = MEM[23846] + MEM[24984];
assign MEM[30091] = MEM[23847] + MEM[26361];
assign MEM[30092] = MEM[23848] + MEM[24544];
assign MEM[30093] = MEM[23849] + MEM[25346];
assign MEM[30094] = MEM[23850] + MEM[28141];
assign MEM[30095] = MEM[23851] + MEM[24194];
assign MEM[30096] = MEM[23852] + MEM[25177];
assign MEM[30097] = MEM[23853] + MEM[24912];
assign MEM[30098] = MEM[23854] + MEM[26291];
assign MEM[30099] = MEM[23855] + MEM[27164];
assign MEM[30100] = MEM[23856] + MEM[24805];
assign MEM[30101] = MEM[23857] + MEM[29331];
assign MEM[30102] = MEM[23858] + MEM[25370];
assign MEM[30103] = MEM[23859] + MEM[26376];
assign MEM[30104] = MEM[23860] + MEM[25274];
assign MEM[30105] = MEM[23861] + MEM[25930];
assign MEM[30106] = MEM[23862] + MEM[24881];
assign MEM[30107] = MEM[23865] + MEM[24908];
assign MEM[30108] = MEM[23866] + MEM[24392];
assign MEM[30109] = MEM[23867] + MEM[26076];
assign MEM[30110] = MEM[23868] + MEM[25316];
assign MEM[30111] = MEM[23869] + MEM[25533];
assign MEM[30112] = MEM[23870] + MEM[24699];
assign MEM[30113] = MEM[23873] + MEM[25407];
assign MEM[30114] = MEM[23874] + MEM[28218];
assign MEM[30115] = MEM[23875] + MEM[28521];
assign MEM[30116] = MEM[23876] + MEM[24309];
assign MEM[30117] = MEM[23877] + MEM[25566];
assign MEM[30118] = MEM[23879] + MEM[24628];
assign MEM[30119] = MEM[23880] + MEM[26321];
assign MEM[30120] = MEM[23881] + MEM[25093];
assign MEM[30121] = MEM[23882] + MEM[25573];
assign MEM[30122] = MEM[23883] + MEM[23951];
assign MEM[30123] = MEM[23884] + MEM[26017];
assign MEM[30124] = MEM[23885] + MEM[26061];
assign MEM[30125] = MEM[23886] + MEM[24749];
assign MEM[30126] = MEM[23887] + MEM[28406];
assign MEM[30127] = MEM[23890] + MEM[25124];
assign MEM[30128] = MEM[23894] + MEM[24842];
assign MEM[30129] = MEM[23895] + MEM[24395];
assign MEM[30130] = MEM[23896] + MEM[26378];
assign MEM[30131] = MEM[23897] + MEM[24476];
assign MEM[30132] = MEM[23898] + MEM[24254];
assign MEM[30133] = MEM[23899] + MEM[27722];
assign MEM[30134] = MEM[23901] + MEM[26913];
assign MEM[30135] = MEM[23903] + MEM[25755];
assign MEM[30136] = MEM[23904] + MEM[28286];
assign MEM[30137] = MEM[23905] + MEM[27791];
assign MEM[30138] = MEM[23906] + MEM[26792];
assign MEM[30139] = MEM[23908] + MEM[24937];
assign MEM[30140] = MEM[23909] + MEM[26927];
assign MEM[30141] = MEM[23910] + MEM[25528];
assign MEM[30142] = MEM[23911] + MEM[28375];
assign MEM[30143] = MEM[23912] + MEM[24454];
assign MEM[30144] = MEM[23913] + MEM[25501];
assign MEM[30145] = MEM[23914] + MEM[25953];
assign MEM[30146] = MEM[23915] + MEM[25100];
assign MEM[30147] = MEM[23916] + MEM[24713];
assign MEM[30148] = MEM[23917] + MEM[25928];
assign MEM[30149] = MEM[23918] + MEM[25014];
assign MEM[30150] = MEM[23919] + MEM[26563];
assign MEM[30151] = MEM[23920] + MEM[25877];
assign MEM[30152] = MEM[23921] + MEM[24610];
assign MEM[30153] = MEM[23923] + MEM[25746];
assign MEM[30154] = MEM[23925] + MEM[24569];
assign MEM[30155] = MEM[23926] + MEM[24589];
assign MEM[30156] = MEM[23927] + MEM[25870];
assign MEM[30157] = MEM[23928] + MEM[24974];
assign MEM[30158] = MEM[23929] + MEM[25602];
assign MEM[30159] = MEM[23931] + MEM[24670];
assign MEM[30160] = MEM[23932] + MEM[26147];
assign MEM[30161] = MEM[23933] + MEM[25086];
assign MEM[30162] = MEM[23934] + MEM[26480];
assign MEM[30163] = MEM[23935] + MEM[26139];
assign MEM[30164] = MEM[23936] + MEM[25944];
assign MEM[30165] = MEM[23937] + MEM[25862];
assign MEM[30166] = MEM[23938] + MEM[23968];
assign MEM[30167] = MEM[23939] + MEM[25459];
assign MEM[30168] = MEM[23941] + MEM[26161];
assign MEM[30169] = MEM[23943] + MEM[25170];
assign MEM[30170] = MEM[23944] + MEM[28913];
assign MEM[30171] = MEM[23945] + MEM[25322];
assign MEM[30172] = MEM[23947] + MEM[26038];
assign MEM[30173] = MEM[23948] + MEM[26787];
assign MEM[30174] = MEM[23949] + MEM[24053];
assign MEM[30175] = MEM[23950] + MEM[25048];
assign MEM[30176] = MEM[23952] + MEM[24350];
assign MEM[30177] = MEM[23953] + MEM[26397];
assign MEM[30178] = MEM[23954] + MEM[25450];
assign MEM[30179] = MEM[23955] + MEM[25373];
assign MEM[30180] = MEM[23956] + MEM[27483];
assign MEM[30181] = MEM[23957] + MEM[24887];
assign MEM[30182] = MEM[23958] + MEM[24882];
assign MEM[30183] = MEM[23959] + MEM[24422];
assign MEM[30184] = MEM[23960] + MEM[27833];
assign MEM[30185] = MEM[23961] + MEM[24752];
assign MEM[30186] = MEM[23962] + MEM[25726];
assign MEM[30187] = MEM[23966] + MEM[26857];
assign MEM[30188] = MEM[23967] + MEM[25493];
assign MEM[30189] = MEM[23969] + MEM[27936];
assign MEM[30190] = MEM[23970] + MEM[27247];
assign MEM[30191] = MEM[23971] + MEM[25175];
assign MEM[30192] = MEM[23973] + MEM[26841];
assign MEM[30193] = MEM[23974] + MEM[25087];
assign MEM[30194] = MEM[23975] + MEM[26552];
assign MEM[30195] = MEM[23976] + MEM[26678];
assign MEM[30196] = MEM[23977] + MEM[25278];
assign MEM[30197] = MEM[23978] + MEM[24547];
assign MEM[30198] = MEM[23980] + MEM[24778];
assign MEM[30199] = MEM[23981] + MEM[25234];
assign MEM[30200] = MEM[23984] + MEM[28074];
assign MEM[30201] = MEM[23986] + MEM[24387];
assign MEM[30202] = MEM[23987] + MEM[25304];
assign MEM[30203] = MEM[23989] + MEM[25590];
assign MEM[30204] = MEM[23990] + MEM[26449];
assign MEM[30205] = MEM[23991] + MEM[28973];
assign MEM[30206] = MEM[23992] + MEM[27471];
assign MEM[30207] = MEM[23993] + MEM[28186];
assign MEM[30208] = MEM[23994] + MEM[27257];
assign MEM[30209] = MEM[23995] + MEM[25122];
assign MEM[30210] = MEM[23996] + MEM[29414];
assign MEM[30211] = MEM[23998] + MEM[26884];
assign MEM[30212] = MEM[23999] + MEM[25624];
assign MEM[30213] = MEM[24000] + MEM[25099];
assign MEM[30214] = MEM[24002] + MEM[26186];
assign MEM[30215] = MEM[24003] + MEM[26045];
assign MEM[30216] = MEM[24006] + MEM[26265];
assign MEM[30217] = MEM[24007] + MEM[25514];
assign MEM[30218] = MEM[24008] + MEM[26183];
assign MEM[30219] = MEM[24009] + MEM[24745];
assign MEM[30220] = MEM[24011] + MEM[29753];
assign MEM[30221] = MEM[24012] + MEM[24382];
assign MEM[30222] = MEM[24014] + MEM[24769];
assign MEM[30223] = MEM[24015] + MEM[28332];
assign MEM[30224] = MEM[24016] + MEM[24884];
assign MEM[30225] = MEM[24017] + MEM[25015];
assign MEM[30226] = MEM[24019] + MEM[25241];
assign MEM[30227] = MEM[24020] + MEM[24592];
assign MEM[30228] = MEM[24021] + MEM[24571];
assign MEM[30229] = MEM[24022] + MEM[26085];
assign MEM[30230] = MEM[24023] + MEM[24259];
assign MEM[30231] = MEM[24031] + MEM[25947];
assign MEM[30232] = MEM[24033] + MEM[24846];
assign MEM[30233] = MEM[24034] + MEM[24920];
assign MEM[30234] = MEM[24035] + MEM[25489];
assign MEM[30235] = MEM[24036] + MEM[27047];
assign MEM[30236] = MEM[24037] + MEM[29012];
assign MEM[30237] = MEM[24038] + MEM[24784];
assign MEM[30238] = MEM[24039] + MEM[27185];
assign MEM[30239] = MEM[24040] + MEM[24883];
assign MEM[30240] = MEM[24041] + MEM[25345];
assign MEM[30241] = MEM[24042] + MEM[26331];
assign MEM[30242] = MEM[24044] + MEM[28584];
assign MEM[30243] = MEM[24045] + MEM[27282];
assign MEM[30244] = MEM[24046] + MEM[25299];
assign MEM[30245] = MEM[24047] + MEM[24838];
assign MEM[30246] = MEM[24048] + MEM[26460];
assign MEM[30247] = MEM[24049] + MEM[25359];
assign MEM[30248] = MEM[24050] + MEM[26467];
assign MEM[30249] = MEM[24051] + MEM[26648];
assign MEM[30250] = MEM[24054] + MEM[26908];
assign MEM[30251] = MEM[24055] + MEM[29178];
assign MEM[30252] = MEM[24056] + MEM[25076];
assign MEM[30253] = MEM[24057] + MEM[25193];
assign MEM[30254] = MEM[24058] + MEM[25654];
assign MEM[30255] = MEM[24059] + MEM[24455];
assign MEM[30256] = MEM[24060] + MEM[26074];
assign MEM[30257] = MEM[24062] + MEM[26535];
assign MEM[30258] = MEM[24063] + MEM[28392];
assign MEM[30259] = MEM[24064] + MEM[26318];
assign MEM[30260] = MEM[24065] + MEM[27544];
assign MEM[30261] = MEM[24066] + MEM[25039];
assign MEM[30262] = MEM[24067] + MEM[24850];
assign MEM[30263] = MEM[24069] + MEM[28730];
assign MEM[30264] = MEM[24070] + MEM[26505];
assign MEM[30265] = MEM[24071] + MEM[24772];
assign MEM[30266] = MEM[24072] + MEM[26121];
assign MEM[30267] = MEM[24073] + MEM[28439];
assign MEM[30268] = MEM[24074] + MEM[24991];
assign MEM[30269] = MEM[24075] + MEM[26078];
assign MEM[30270] = MEM[24076] + MEM[27542];
assign MEM[30271] = MEM[24077] + MEM[29458];
assign MEM[30272] = MEM[24079] + MEM[26313];
assign MEM[30273] = MEM[24080] + MEM[24310];
assign MEM[30274] = MEM[24081] + MEM[25655];
assign MEM[30275] = MEM[24083] + MEM[25464];
assign MEM[30276] = MEM[24084] + MEM[27195];
assign MEM[30277] = MEM[24087] + MEM[25567];
assign MEM[30278] = MEM[24088] + MEM[26191];
assign MEM[30279] = MEM[24089] + MEM[28487];
assign MEM[30280] = MEM[24090] + MEM[25789];
assign MEM[30281] = MEM[24091] + MEM[27352];
assign MEM[30282] = MEM[24092] + MEM[25102];
assign MEM[30283] = MEM[24093] + MEM[26355];
assign MEM[30284] = MEM[24094] + MEM[27226];
assign MEM[30285] = MEM[24096] + MEM[25136];
assign MEM[30286] = MEM[24098] + MEM[25440];
assign MEM[30287] = MEM[24100] + MEM[24896];
assign MEM[30288] = MEM[24101] + MEM[26225];
assign MEM[30289] = MEM[24102] + MEM[26266];
assign MEM[30290] = MEM[24103] + MEM[26022];
assign MEM[30291] = MEM[24104] + MEM[25535];
assign MEM[30292] = MEM[24105] + MEM[25684];
assign MEM[30293] = MEM[24106] + MEM[24933];
assign MEM[30294] = MEM[24108] + MEM[28930];
assign MEM[30295] = MEM[24109] + MEM[24728];
assign MEM[30296] = MEM[24110] + MEM[26888];
assign MEM[30297] = MEM[24111] + MEM[25673];
assign MEM[30298] = MEM[24112] + MEM[26718];
assign MEM[30299] = MEM[24113] + MEM[27981];
assign MEM[30300] = MEM[24115] + MEM[24847];
assign MEM[30301] = MEM[24117] + MEM[28743];
assign MEM[30302] = MEM[24118] + MEM[24142];
assign MEM[30303] = MEM[24119] + MEM[24602];
assign MEM[30304] = MEM[24121] + MEM[28073];
assign MEM[30305] = MEM[24123] + MEM[26504];
assign MEM[30306] = MEM[24126] + MEM[28818];
assign MEM[30307] = MEM[24127] + MEM[25851];
assign MEM[30308] = MEM[24128] + MEM[25596];
assign MEM[30309] = MEM[24129] + MEM[25751];
assign MEM[30310] = MEM[24130] + MEM[26915];
assign MEM[30311] = MEM[24131] + MEM[26860];
assign MEM[30312] = MEM[24132] + MEM[26215];
assign MEM[30313] = MEM[24133] + MEM[26941];
assign MEM[30314] = MEM[24134] + MEM[24389];
assign MEM[30315] = MEM[24135] + MEM[26854];
assign MEM[30316] = MEM[24136] + MEM[25592];
assign MEM[30317] = MEM[24137] + MEM[27996];
assign MEM[30318] = MEM[24138] + MEM[24746];
assign MEM[30319] = MEM[24139] + MEM[25405];
assign MEM[30320] = MEM[24140] + MEM[24542];
assign MEM[30321] = MEM[24141] + MEM[25912];
assign MEM[30322] = MEM[24143] + MEM[28028];
assign MEM[30323] = MEM[24144] + MEM[24539];
assign MEM[30324] = MEM[24145] + MEM[24844];
assign MEM[30325] = MEM[24147] + MEM[26624];
assign MEM[30326] = MEM[24148] + MEM[27200];
assign MEM[30327] = MEM[24149] + MEM[27028];
assign MEM[30328] = MEM[24151] + MEM[25557];
assign MEM[30329] = MEM[24152] + MEM[25882];
assign MEM[30330] = MEM[24154] + MEM[24341];
assign MEM[30331] = MEM[24155] + MEM[27605];
assign MEM[30332] = MEM[24156] + MEM[24580];
assign MEM[30333] = MEM[24157] + MEM[26577];
assign MEM[30334] = MEM[24158] + MEM[26481];
assign MEM[30335] = MEM[24159] + MEM[26815];
assign MEM[30336] = MEM[24161] + MEM[26184];
assign MEM[30337] = MEM[24163] + MEM[25394];
assign MEM[30338] = MEM[24164] + MEM[29239];
assign MEM[30339] = MEM[24165] + MEM[26767];
assign MEM[30340] = MEM[24168] + MEM[24509];
assign MEM[30341] = MEM[24169] + MEM[25239];
assign MEM[30342] = MEM[24170] + MEM[24986];
assign MEM[30343] = MEM[24171] + MEM[26532];
assign MEM[30344] = MEM[24172] + MEM[26033];
assign MEM[30345] = MEM[24174] + MEM[24690];
assign MEM[30346] = MEM[24175] + MEM[26468];
assign MEM[30347] = MEM[24176] + MEM[25472];
assign MEM[30348] = MEM[24177] + MEM[26229];
assign MEM[30349] = MEM[24178] + MEM[24989];
assign MEM[30350] = MEM[24182] + MEM[25515];
assign MEM[30351] = MEM[24183] + MEM[27988];
assign MEM[30352] = MEM[24184] + MEM[26962];
assign MEM[30353] = MEM[24185] + MEM[26905];
assign MEM[30354] = MEM[24187] + MEM[25706];
assign MEM[30355] = MEM[24188] + MEM[26725];
assign MEM[30356] = MEM[24190] + MEM[25729];
assign MEM[30357] = MEM[24191] + MEM[26510];
assign MEM[30358] = MEM[24192] + MEM[24687];
assign MEM[30359] = MEM[24193] + MEM[26350];
assign MEM[30360] = MEM[24195] + MEM[26129];
assign MEM[30361] = MEM[24196] + MEM[27386];
assign MEM[30362] = MEM[24197] + MEM[24970];
assign MEM[30363] = MEM[24199] + MEM[26591];
assign MEM[30364] = MEM[24200] + MEM[26448];
assign MEM[30365] = MEM[24201] + MEM[24757];
assign MEM[30366] = MEM[24205] + MEM[26010];
assign MEM[30367] = MEM[24206] + MEM[24435];
assign MEM[30368] = MEM[24207] + MEM[29028];
assign MEM[30369] = MEM[24209] + MEM[24737];
assign MEM[30370] = MEM[24210] + MEM[24999];
assign MEM[30371] = MEM[24213] + MEM[24267];
assign MEM[30372] = MEM[24214] + MEM[25992];
assign MEM[30373] = MEM[24215] + MEM[26206];
assign MEM[30374] = MEM[24216] + MEM[26593];
assign MEM[30375] = MEM[24217] + MEM[25509];
assign MEM[30376] = MEM[24219] + MEM[27531];
assign MEM[30377] = MEM[24220] + MEM[26011];
assign MEM[30378] = MEM[24222] + MEM[26185];
assign MEM[30379] = MEM[24224] + MEM[25932];
assign MEM[30380] = MEM[24225] + MEM[26404];
assign MEM[30381] = MEM[24226] + MEM[25665];
assign MEM[30382] = MEM[24227] + MEM[26471];
assign MEM[30383] = MEM[24228] + MEM[26120];
assign MEM[30384] = MEM[24229] + MEM[25194];
assign MEM[30385] = MEM[24230] + MEM[26131];
assign MEM[30386] = MEM[24231] + MEM[26243];
assign MEM[30387] = MEM[24233] + MEM[27217];
assign MEM[30388] = MEM[24234] + MEM[25313];
assign MEM[30389] = MEM[24235] + MEM[27954];
assign MEM[30390] = MEM[24236] + MEM[26619];
assign MEM[30391] = MEM[24237] + MEM[25222];
assign MEM[30392] = MEM[24239] + MEM[26626];
assign MEM[30393] = MEM[24240] + MEM[27100];
assign MEM[30394] = MEM[24241] + MEM[26509];
assign MEM[30395] = MEM[24242] + MEM[25457];
assign MEM[30396] = MEM[24243] + MEM[24513];
assign MEM[30397] = MEM[24244] + MEM[25041];
assign MEM[30398] = MEM[24245] + MEM[25707];
assign MEM[30399] = MEM[24246] + MEM[25310];
assign MEM[30400] = MEM[24247] + MEM[25815];
assign MEM[30401] = MEM[24248] + MEM[27776];
assign MEM[30402] = MEM[24249] + MEM[25071];
assign MEM[30403] = MEM[24250] + MEM[25942];
assign MEM[30404] = MEM[24251] + MEM[27410];
assign MEM[30405] = MEM[24252] + MEM[25326];
assign MEM[30406] = MEM[24253] + MEM[27054];
assign MEM[30407] = MEM[24255] + MEM[25583];
assign MEM[30408] = MEM[24256] + MEM[26955];
assign MEM[30409] = MEM[24257] + MEM[25772];
assign MEM[30410] = MEM[24258] + MEM[26729];
assign MEM[30411] = MEM[24260] + MEM[25641];
assign MEM[30412] = MEM[24261] + MEM[25258];
assign MEM[30413] = MEM[24262] + MEM[26720];
assign MEM[30414] = MEM[24263] + MEM[26219];
assign MEM[30415] = MEM[24264] + MEM[25438];
assign MEM[30416] = MEM[24265] + MEM[26979];
assign MEM[30417] = MEM[24266] + MEM[25189];
assign MEM[30418] = MEM[24269] + MEM[26261];
assign MEM[30419] = MEM[24270] + MEM[28037];
assign MEM[30420] = MEM[24271] + MEM[26371];
assign MEM[30421] = MEM[24272] + MEM[26388];
assign MEM[30422] = MEM[24273] + MEM[26255];
assign MEM[30423] = MEM[24274] + MEM[27066];
assign MEM[30424] = MEM[24275] + MEM[25891];
assign MEM[30425] = MEM[24276] + MEM[25393];
assign MEM[30426] = MEM[24278] + MEM[25696];
assign MEM[30427] = MEM[24279] + MEM[26268];
assign MEM[30428] = MEM[24281] + MEM[24545];
assign MEM[30429] = MEM[24282] + MEM[25820];
assign MEM[30430] = MEM[24284] + MEM[26896];
assign MEM[30431] = MEM[24285] + MEM[24928];
assign MEM[30432] = MEM[24287] + MEM[26278];
assign MEM[30433] = MEM[24288] + MEM[26068];
assign MEM[30434] = MEM[24289] + MEM[26375];
assign MEM[30435] = MEM[24291] + MEM[24819];
assign MEM[30436] = MEM[24292] + MEM[26124];
assign MEM[30437] = MEM[24293] + MEM[25587];
assign MEM[30438] = MEM[24294] + MEM[27736];
assign MEM[30439] = MEM[24295] + MEM[25925];
assign MEM[30440] = MEM[24300] + MEM[24825];
assign MEM[30441] = MEM[24301] + MEM[25988];
assign MEM[30442] = MEM[24302] + MEM[26242];
assign MEM[30443] = MEM[24303] + MEM[26230];
assign MEM[30444] = MEM[24304] + MEM[27317];
assign MEM[30445] = MEM[24305] + MEM[24565];
assign MEM[30446] = MEM[24306] + MEM[25970];
assign MEM[30447] = MEM[24308] + MEM[26381];
assign MEM[30448] = MEM[24311] + MEM[25290];
assign MEM[30449] = MEM[24312] + MEM[25698];
assign MEM[30450] = MEM[24313] + MEM[25761];
assign MEM[30451] = MEM[24314] + MEM[25685];
assign MEM[30452] = MEM[24315] + MEM[25259];
assign MEM[30453] = MEM[24316] + MEM[26253];
assign MEM[30454] = MEM[24318] + MEM[25251];
assign MEM[30455] = MEM[24319] + MEM[25031];
assign MEM[30456] = MEM[24320] + MEM[25734];
assign MEM[30457] = MEM[24322] + MEM[28292];
assign MEM[30458] = MEM[24324] + MEM[25279];
assign MEM[30459] = MEM[24325] + MEM[26037];
assign MEM[30460] = MEM[24326] + MEM[24812];
assign MEM[30461] = MEM[24327] + MEM[26167];
assign MEM[30462] = MEM[24330] + MEM[26394];
assign MEM[30463] = MEM[24331] + MEM[25739];
assign MEM[30464] = MEM[24332] + MEM[25672];
assign MEM[30465] = MEM[24334] + MEM[25804];
assign MEM[30466] = MEM[24337] + MEM[24674];
assign MEM[30467] = MEM[24338] + MEM[26001];
assign MEM[30468] = MEM[24339] + MEM[28965];
assign MEM[30469] = MEM[24340] + MEM[25786];
assign MEM[30470] = MEM[24342] + MEM[25517];
assign MEM[30471] = MEM[24343] + MEM[28116];
assign MEM[30472] = MEM[24344] + MEM[25069];
assign MEM[30473] = MEM[24345] + MEM[26007];
assign MEM[30474] = MEM[24346] + MEM[25433];
assign MEM[30475] = MEM[24347] + MEM[25554];
assign MEM[30476] = MEM[24348] + MEM[26662];
assign MEM[30477] = MEM[24351] + MEM[25878];
assign MEM[30478] = MEM[24352] + MEM[25807];
assign MEM[30479] = MEM[24354] + MEM[25208];
assign MEM[30480] = MEM[24355] + MEM[27396];
assign MEM[30481] = MEM[24358] + MEM[25430];
assign MEM[30482] = MEM[24360] + MEM[26588];
assign MEM[30483] = MEM[24361] + MEM[25917];
assign MEM[30484] = MEM[24362] + MEM[25337];
assign MEM[30485] = MEM[24363] + MEM[25968];
assign MEM[30486] = MEM[24365] + MEM[26649];
assign MEM[30487] = MEM[24366] + MEM[25281];
assign MEM[30488] = MEM[24367] + MEM[26549];
assign MEM[30489] = MEM[24368] + MEM[26352];
assign MEM[30490] = MEM[24369] + MEM[25598];
assign MEM[30491] = MEM[24371] + MEM[25883];
assign MEM[30492] = MEM[24372] + MEM[25180];
assign MEM[30493] = MEM[24373] + MEM[25496];
assign MEM[30494] = MEM[24375] + MEM[28690];
assign MEM[30495] = MEM[24376] + MEM[25771];
assign MEM[30496] = MEM[24377] + MEM[26351];
assign MEM[30497] = MEM[24378] + MEM[26041];
assign MEM[30498] = MEM[24380] + MEM[27401];
assign MEM[30499] = MEM[24381] + MEM[27076];
assign MEM[30500] = MEM[24383] + MEM[26646];
assign MEM[30501] = MEM[24384] + MEM[25785];
assign MEM[30502] = MEM[24385] + MEM[25788];
assign MEM[30503] = MEM[24388] + MEM[26922];
assign MEM[30504] = MEM[24390] + MEM[26240];
assign MEM[30505] = MEM[24393] + MEM[26553];
assign MEM[30506] = MEM[24396] + MEM[25495];
assign MEM[30507] = MEM[24397] + MEM[26281];
assign MEM[30508] = MEM[24398] + MEM[25399];
assign MEM[30509] = MEM[24399] + MEM[27005];
assign MEM[30510] = MEM[24401] + MEM[24863];
assign MEM[30511] = MEM[24402] + MEM[25130];
assign MEM[30512] = MEM[24403] + MEM[25132];
assign MEM[30513] = MEM[24404] + MEM[25542];
assign MEM[30514] = MEM[24405] + MEM[25118];
assign MEM[30515] = MEM[24406] + MEM[28794];
assign MEM[30516] = MEM[24407] + MEM[26807];
assign MEM[30517] = MEM[24410] + MEM[27287];
assign MEM[30518] = MEM[24411] + MEM[26782];
assign MEM[30519] = MEM[24412] + MEM[26617];
assign MEM[30520] = MEM[24413] + MEM[25893];
assign MEM[30521] = MEM[24414] + MEM[24787];
assign MEM[30522] = MEM[24415] + MEM[24663];
assign MEM[30523] = MEM[24416] + MEM[25683];
assign MEM[30524] = MEM[24417] + MEM[25984];
assign MEM[30525] = MEM[24418] + MEM[27221];
assign MEM[30526] = MEM[24419] + MEM[27620];
assign MEM[30527] = MEM[24420] + MEM[25188];
assign MEM[30528] = MEM[24421] + MEM[26105];
assign MEM[30529] = MEM[24423] + MEM[25420];
assign MEM[30530] = MEM[24424] + MEM[24709];
assign MEM[30531] = MEM[24427] + MEM[25417];
assign MEM[30532] = MEM[24428] + MEM[25794];
assign MEM[30533] = MEM[24429] + MEM[25458];
assign MEM[30534] = MEM[24430] + MEM[28418];
assign MEM[30535] = MEM[24431] + MEM[26682];
assign MEM[30536] = MEM[24432] + MEM[25138];
assign MEM[30537] = MEM[24434] + MEM[25519];
assign MEM[30538] = MEM[24436] + MEM[26902];
assign MEM[30539] = MEM[24437] + MEM[25174];
assign MEM[30540] = MEM[24440] + MEM[25671];
assign MEM[30541] = MEM[24442] + MEM[26578];
assign MEM[30542] = MEM[24443] + MEM[24973];
assign MEM[30543] = MEM[24444] + MEM[25023];
assign MEM[30544] = MEM[24445] + MEM[26683];
assign MEM[30545] = MEM[24446] + MEM[26486];
assign MEM[30546] = MEM[24450] + MEM[25619];
assign MEM[30547] = MEM[24452] + MEM[26058];
assign MEM[30548] = MEM[24453] + MEM[27371];
assign MEM[30549] = MEM[24456] + MEM[26607];
assign MEM[30550] = MEM[24457] + MEM[28735];
assign MEM[30551] = MEM[24458] + MEM[27417];
assign MEM[30552] = MEM[24459] + MEM[26250];
assign MEM[30553] = MEM[24462] + MEM[27792];
assign MEM[30554] = MEM[24463] + MEM[27914];
assign MEM[30555] = MEM[24465] + MEM[28065];
assign MEM[30556] = MEM[24466] + MEM[25996];
assign MEM[30557] = MEM[24467] + MEM[26027];
assign MEM[30558] = MEM[24468] + MEM[25599];
assign MEM[30559] = MEM[24470] + MEM[26358];
assign MEM[30560] = MEM[24471] + MEM[25488];
assign MEM[30561] = MEM[24472] + MEM[24826];
assign MEM[30562] = MEM[24473] + MEM[26288];
assign MEM[30563] = MEM[24474] + MEM[24915];
assign MEM[30564] = MEM[24475] + MEM[26132];
assign MEM[30565] = MEM[24477] + MEM[25277];
assign MEM[30566] = MEM[24478] + MEM[28762];
assign MEM[30567] = MEM[24479] + MEM[25314];
assign MEM[30568] = MEM[24480] + MEM[27985];
assign MEM[30569] = MEM[24482] + MEM[25833];
assign MEM[30570] = MEM[24483] + MEM[25143];
assign MEM[30571] = MEM[24484] + MEM[25406];
assign MEM[30572] = MEM[24486] + MEM[24824];
assign MEM[30573] = MEM[24488] + MEM[25034];
assign MEM[30574] = MEM[24489] + MEM[27344];
assign MEM[30575] = MEM[24490] + MEM[26320];
assign MEM[30576] = MEM[24491] + MEM[25889];
assign MEM[30577] = MEM[24492] + MEM[24935];
assign MEM[30578] = MEM[24493] + MEM[25896];
assign MEM[30579] = MEM[24494] + MEM[25007];
assign MEM[30580] = MEM[24495] + MEM[28350];
assign MEM[30581] = MEM[24496] + MEM[28047];
assign MEM[30582] = MEM[24499] + MEM[25594];
assign MEM[30583] = MEM[24500] + MEM[25141];
assign MEM[30584] = MEM[24501] + MEM[25368];
assign MEM[30585] = MEM[24502] + MEM[26067];
assign MEM[30586] = MEM[24503] + MEM[29021];
assign MEM[30587] = MEM[24504] + MEM[27263];
assign MEM[30588] = MEM[24506] + MEM[26403];
assign MEM[30589] = MEM[24507] + MEM[27090];
assign MEM[30590] = MEM[24512] + MEM[24828];
assign MEM[30591] = MEM[24515] + MEM[25101];
assign MEM[30592] = MEM[24516] + MEM[26116];
assign MEM[30593] = MEM[24517] + MEM[25161];
assign MEM[30594] = MEM[24518] + MEM[26930];
assign MEM[30595] = MEM[24519] + MEM[28136];
assign MEM[30596] = MEM[24520] + MEM[25895];
assign MEM[30597] = MEM[24522] + MEM[25916];
assign MEM[30598] = MEM[24525] + MEM[26759];
assign MEM[30599] = MEM[24526] + MEM[26983];
assign MEM[30600] = MEM[24527] + MEM[26008];
assign MEM[30601] = MEM[24528] + MEM[29685];
assign MEM[30602] = MEM[24530] + MEM[25167];
assign MEM[30603] = MEM[24531] + MEM[27058];
assign MEM[30604] = MEM[24532] + MEM[25283];
assign MEM[30605] = MEM[24533] + MEM[24917];
assign MEM[30606] = MEM[24535] + MEM[28853];
assign MEM[30607] = MEM[24536] + MEM[25666];
assign MEM[30608] = MEM[24537] + MEM[25579];
assign MEM[30609] = MEM[24538] + MEM[24742];
assign MEM[30610] = MEM[24541] + MEM[27658];
assign MEM[30611] = MEM[24543] + MEM[26919];
assign MEM[30612] = MEM[24546] + MEM[26494];
assign MEM[30613] = MEM[24548] + MEM[28776];
assign MEM[30614] = MEM[24549] + MEM[27582];
assign MEM[30615] = MEM[24550] + MEM[24586];
assign MEM[30616] = MEM[24553] + MEM[24880];
assign MEM[30617] = MEM[24554] + MEM[27422];
assign MEM[30618] = MEM[24556] + MEM[27541];
assign MEM[30619] = MEM[24558] + MEM[28077];
assign MEM[30620] = MEM[24560] + MEM[29125];
assign MEM[30621] = MEM[24561] + MEM[26195];
assign MEM[30622] = MEM[24562] + MEM[27557];
assign MEM[30623] = MEM[24563] + MEM[28321];
assign MEM[30624] = MEM[24567] + MEM[25728];
assign MEM[30625] = MEM[24568] + MEM[28959];
assign MEM[30626] = MEM[24570] + MEM[26688];
assign MEM[30627] = MEM[24572] + MEM[25875];
assign MEM[30628] = MEM[24573] + MEM[27598];
assign MEM[30629] = MEM[24575] + MEM[26575];
assign MEM[30630] = MEM[24576] + MEM[27360];
assign MEM[30631] = MEM[24577] + MEM[25197];
assign MEM[30632] = MEM[24578] + MEM[27072];
assign MEM[30633] = MEM[24579] + MEM[25898];
assign MEM[30634] = MEM[24581] + MEM[24801];
assign MEM[30635] = MEM[24582] + MEM[29023];
assign MEM[30636] = MEM[24583] + MEM[27278];
assign MEM[30637] = MEM[24584] + MEM[26316];
assign MEM[30638] = MEM[24585] + MEM[25461];
assign MEM[30639] = MEM[24588] + MEM[25808];
assign MEM[30640] = MEM[24590] + MEM[28050];
assign MEM[30641] = MEM[24593] + MEM[26337];
assign MEM[30642] = MEM[24595] + MEM[26802];
assign MEM[30643] = MEM[24596] + MEM[27349];
assign MEM[30644] = MEM[24598] + MEM[26286];
assign MEM[30645] = MEM[24599] + MEM[26880];
assign MEM[30646] = MEM[24601] + MEM[25228];
assign MEM[30647] = MEM[24603] + MEM[26140];
assign MEM[30648] = MEM[24604] + MEM[25155];
assign MEM[30649] = MEM[24606] + MEM[25376];
assign MEM[30650] = MEM[24607] + MEM[25383];
assign MEM[30651] = MEM[24608] + MEM[25042];
assign MEM[30652] = MEM[24613] + MEM[25563];
assign MEM[30653] = MEM[24614] + MEM[26707];
assign MEM[30654] = MEM[24615] + MEM[25253];
assign MEM[30655] = MEM[24616] + MEM[26249];
assign MEM[30656] = MEM[24617] + MEM[27440];
assign MEM[30657] = MEM[24618] + MEM[26485];
assign MEM[30658] = MEM[24620] + MEM[24916];
assign MEM[30659] = MEM[24621] + MEM[25888];
assign MEM[30660] = MEM[24622] + MEM[25227];
assign MEM[30661] = MEM[24625] + MEM[28790];
assign MEM[30662] = MEM[24626] + MEM[25271];
assign MEM[30663] = MEM[24627] + MEM[25543];
assign MEM[30664] = MEM[24629] + MEM[27870];
assign MEM[30665] = MEM[24630] + MEM[25718];
assign MEM[30666] = MEM[24632] + MEM[24848];
assign MEM[30667] = MEM[24633] + MEM[26497];
assign MEM[30668] = MEM[24634] + MEM[25152];
assign MEM[30669] = MEM[24636] + MEM[26452];
assign MEM[30670] = MEM[24638] + MEM[26751];
assign MEM[30671] = MEM[24639] + MEM[27149];
assign MEM[30672] = MEM[24640] + MEM[25486];
assign MEM[30673] = MEM[24642] + MEM[26149];
assign MEM[30674] = MEM[24645] + MEM[28754];
assign MEM[30675] = MEM[24646] + MEM[25622];
assign MEM[30676] = MEM[24648] + MEM[26168];
assign MEM[30677] = MEM[24649] + MEM[25302];
assign MEM[30678] = MEM[24650] + MEM[25004];
assign MEM[30679] = MEM[24651] + MEM[26818];
assign MEM[30680] = MEM[24653] + MEM[25873];
assign MEM[30681] = MEM[24655] + MEM[25544];
assign MEM[30682] = MEM[24657] + MEM[27563];
assign MEM[30683] = MEM[24658] + MEM[26342];
assign MEM[30684] = MEM[24659] + MEM[24776];
assign MEM[30685] = MEM[24660] + MEM[25679];
assign MEM[30686] = MEM[24661] + MEM[29228];
assign MEM[30687] = MEM[24662] + MEM[25959];
assign MEM[30688] = MEM[24664] + MEM[26727];
assign MEM[30689] = MEM[24665] + MEM[26256];
assign MEM[30690] = MEM[24666] + MEM[24953];
assign MEM[30691] = MEM[24668] + MEM[25478];
assign MEM[30692] = MEM[24669] + MEM[25291];
assign MEM[30693] = MEM[24671] + MEM[26566];
assign MEM[30694] = MEM[24672] + MEM[25315];
assign MEM[30695] = MEM[24673] + MEM[28545];
assign MEM[30696] = MEM[24675] + MEM[26760];
assign MEM[30697] = MEM[24676] + MEM[28256];
assign MEM[30698] = MEM[24679] + MEM[28635];
assign MEM[30699] = MEM[24681] + MEM[27250];
assign MEM[30700] = MEM[24682] + MEM[25871];
assign MEM[30701] = MEM[24683] + MEM[26918];
assign MEM[30702] = MEM[24684] + MEM[27719];
assign MEM[30703] = MEM[24688] + MEM[25358];
assign MEM[30704] = MEM[24689] + MEM[26805];
assign MEM[30705] = MEM[24691] + MEM[26095];
assign MEM[30706] = MEM[24692] + MEM[26379];
assign MEM[30707] = MEM[24693] + MEM[25200];
assign MEM[30708] = MEM[24696] + MEM[26329];
assign MEM[30709] = MEM[24698] + MEM[25173];
assign MEM[30710] = MEM[24701] + MEM[25319];
assign MEM[30711] = MEM[24702] + MEM[26164];
assign MEM[30712] = MEM[24703] + MEM[28326];
assign MEM[30713] = MEM[24704] + MEM[25073];
assign MEM[30714] = MEM[24705] + MEM[25425];
assign MEM[30715] = MEM[24706] + MEM[26442];
assign MEM[30716] = MEM[24707] + MEM[26495];
assign MEM[30717] = MEM[24708] + MEM[25360];
assign MEM[30718] = MEM[24710] + MEM[27656];
assign MEM[30719] = MEM[24711] + MEM[27262];
assign MEM[30720] = MEM[24714] + MEM[26900];
assign MEM[30721] = MEM[24715] + MEM[25166];
assign MEM[30722] = MEM[24716] + MEM[28624];
assign MEM[30723] = MEM[24719] + MEM[26706];
assign MEM[30724] = MEM[24720] + MEM[26812];
assign MEM[30725] = MEM[24721] + MEM[28459];
assign MEM[30726] = MEM[24722] + MEM[26711];
assign MEM[30727] = MEM[24723] + MEM[25580];
assign MEM[30728] = MEM[24724] + MEM[25400];
assign MEM[30729] = MEM[24725] + MEM[26881];
assign MEM[30730] = MEM[24726] + MEM[25513];
assign MEM[30731] = MEM[24727] + MEM[27881];
assign MEM[30732] = MEM[24730] + MEM[28181];
assign MEM[30733] = MEM[24731] + MEM[28989];
assign MEM[30734] = MEM[24732] + MEM[25843];
assign MEM[30735] = MEM[24735] + MEM[25950];
assign MEM[30736] = MEM[24736] + MEM[26541];
assign MEM[30737] = MEM[24739] + MEM[25018];
assign MEM[30738] = MEM[24740] + MEM[27150];
assign MEM[30739] = MEM[24743] + MEM[25182];
assign MEM[30740] = MEM[24748] + MEM[25038];
assign MEM[30741] = MEM[24751] + MEM[25644];
assign MEM[30742] = MEM[24753] + MEM[24865];
assign MEM[30743] = MEM[24754] + MEM[25850];
assign MEM[30744] = MEM[24755] + MEM[25043];
assign MEM[30745] = MEM[24759] + MEM[28758];
assign MEM[30746] = MEM[24760] + MEM[26317];
assign MEM[30747] = MEM[24762] + MEM[26146];
assign MEM[30748] = MEM[24763] + MEM[25687];
assign MEM[30749] = MEM[24764] + MEM[26730];
assign MEM[30750] = MEM[24765] + MEM[26112];
assign MEM[30751] = MEM[24766] + MEM[28154];
assign MEM[30752] = MEM[24767] + MEM[26025];
assign MEM[30753] = MEM[24768] + MEM[26784];
assign MEM[30754] = MEM[24770] + MEM[27521];
assign MEM[30755] = MEM[24771] + MEM[25331];
assign MEM[30756] = MEM[24773] + MEM[24936];
assign MEM[30757] = MEM[24774] + MEM[26006];
assign MEM[30758] = MEM[24775] + MEM[26441];
assign MEM[30759] = MEM[24777] + MEM[25694];
assign MEM[30760] = MEM[24779] + MEM[29381];
assign MEM[30761] = MEM[24781] + MEM[28026];
assign MEM[30762] = MEM[24783] + MEM[26165];
assign MEM[30763] = MEM[24786] + MEM[26929];
assign MEM[30764] = MEM[24789] + MEM[26203];
assign MEM[30765] = MEM[24791] + MEM[25651];
assign MEM[30766] = MEM[24792] + MEM[25939];
assign MEM[30767] = MEM[24793] + MEM[25199];
assign MEM[30768] = MEM[24794] + MEM[26597];
assign MEM[30769] = MEM[24796] + MEM[28975];
assign MEM[30770] = MEM[24798] + MEM[29439];
assign MEM[30771] = MEM[24799] + MEM[25057];
assign MEM[30772] = MEM[24800] + MEM[25633];
assign MEM[30773] = MEM[24802] + MEM[27896];
assign MEM[30774] = MEM[24803] + MEM[27248];
assign MEM[30775] = MEM[24804] + MEM[25980];
assign MEM[30776] = MEM[24806] + MEM[29734];
assign MEM[30777] = MEM[24808] + MEM[26762];
assign MEM[30778] = MEM[24810] + MEM[28520];
assign MEM[30779] = MEM[24811] + MEM[26651];
assign MEM[30780] = MEM[24816] + MEM[25108];
assign MEM[30781] = MEM[24817] + MEM[25190];
assign MEM[30782] = MEM[24818] + MEM[25202];
assign MEM[30783] = MEM[24821] + MEM[28373];
assign MEM[30784] = MEM[24822] + MEM[28243];
assign MEM[30785] = MEM[24827] + MEM[25408];
assign MEM[30786] = MEM[24829] + MEM[25432];
assign MEM[30787] = MEM[24831] + MEM[28129];
assign MEM[30788] = MEM[24833] + MEM[28083];
assign MEM[30789] = MEM[24834] + MEM[29243];
assign MEM[30790] = MEM[24835] + MEM[26435];
assign MEM[30791] = MEM[24836] + MEM[26145];
assign MEM[30792] = MEM[24837] + MEM[26621];
assign MEM[30793] = MEM[24839] + MEM[25803];
assign MEM[30794] = MEM[24840] + MEM[25565];
assign MEM[30795] = MEM[24854] + MEM[25492];
assign MEM[30796] = MEM[24855] + MEM[25483];
assign MEM[30797] = MEM[24856] + MEM[28189];
assign MEM[30798] = MEM[24857] + MEM[27728];
assign MEM[30799] = MEM[24858] + MEM[27664];
assign MEM[30800] = MEM[24859] + MEM[26142];
assign MEM[30801] = MEM[24861] + MEM[25921];
assign MEM[30802] = MEM[24862] + MEM[26455];
assign MEM[30803] = MEM[24864] + MEM[26334];
assign MEM[30804] = MEM[24866] + MEM[26392];
assign MEM[30805] = MEM[24869] + MEM[24971];
assign MEM[30806] = MEM[24871] + MEM[25377];
assign MEM[30807] = MEM[24873] + MEM[27351];
assign MEM[30808] = MEM[24874] + MEM[25353];
assign MEM[30809] = MEM[24876] + MEM[26436];
assign MEM[30810] = MEM[24877] + MEM[27980];
assign MEM[30811] = MEM[24878] + MEM[25421];
assign MEM[30812] = MEM[24879] + MEM[27038];
assign MEM[30813] = MEM[24885] + MEM[25568];
assign MEM[30814] = MEM[24886] + MEM[27420];
assign MEM[30815] = MEM[24888] + MEM[26750];
assign MEM[30816] = MEM[24889] + MEM[26712];
assign MEM[30817] = MEM[24890] + MEM[25708];
assign MEM[30818] = MEM[24894] + MEM[25886];
assign MEM[30819] = MEM[24895] + MEM[25191];
assign MEM[30820] = MEM[24898] + MEM[27031];
assign MEM[30821] = MEM[24899] + MEM[26108];
assign MEM[30822] = MEM[24901] + MEM[26659];
assign MEM[30823] = MEM[24902] + MEM[25692];
assign MEM[30824] = MEM[24903] + MEM[28274];
assign MEM[30825] = MEM[24904] + MEM[26415];
assign MEM[30826] = MEM[24905] + MEM[28662];
assign MEM[30827] = MEM[24906] + MEM[27597];
assign MEM[30828] = MEM[24907] + MEM[26285];
assign MEM[30829] = MEM[24909] + MEM[26372];
assign MEM[30830] = MEM[24911] + MEM[25773];
assign MEM[30831] = MEM[24913] + MEM[25225];
assign MEM[30832] = MEM[24919] + MEM[25720];
assign MEM[30833] = MEM[24922] + MEM[26744];
assign MEM[30834] = MEM[24923] + MEM[26890];
assign MEM[30835] = MEM[24924] + MEM[26263];
assign MEM[30836] = MEM[24926] + MEM[27279];
assign MEM[30837] = MEM[24927] + MEM[25691];
assign MEM[30838] = MEM[24929] + MEM[25775];
assign MEM[30839] = MEM[24930] + MEM[25662];
assign MEM[30840] = MEM[24931] + MEM[26465];
assign MEM[30841] = MEM[24932] + MEM[26075];
assign MEM[30842] = MEM[24934] + MEM[26570];
assign MEM[30843] = MEM[24938] + MEM[26133];
assign MEM[30844] = MEM[24939] + MEM[25607];
assign MEM[30845] = MEM[24941] + MEM[25419];
assign MEM[30846] = MEM[24942] + MEM[27346];
assign MEM[30847] = MEM[24945] + MEM[26833];
assign MEM[30848] = MEM[24946] + MEM[25818];
assign MEM[30849] = MEM[24947] + MEM[26042];
assign MEM[30850] = MEM[24949] + MEM[25682];
assign MEM[30851] = MEM[24950] + MEM[25806];
assign MEM[30852] = MEM[24951] + MEM[28560];
assign MEM[30853] = MEM[24952] + MEM[25094];
assign MEM[30854] = MEM[24954] + MEM[25550];
assign MEM[30855] = MEM[24955] + MEM[26373];
assign MEM[30856] = MEM[24956] + MEM[29497];
assign MEM[30857] = MEM[24959] + MEM[26852];
assign MEM[30858] = MEM[24960] + MEM[27394];
assign MEM[30859] = MEM[24961] + MEM[27337];
assign MEM[30860] = MEM[24962] + MEM[26489];
assign MEM[30861] = MEM[24963] + MEM[25540];
assign MEM[30862] = MEM[24965] + MEM[25774];
assign MEM[30863] = MEM[24967] + MEM[27171];
assign MEM[30864] = MEM[24969] + MEM[25936];
assign MEM[30865] = MEM[24972] + MEM[25948];
assign MEM[30866] = MEM[24975] + MEM[26778];
assign MEM[30867] = MEM[24977] + MEM[25287];
assign MEM[30868] = MEM[24978] + MEM[25525];
assign MEM[30869] = MEM[24979] + MEM[25961];
assign MEM[30870] = MEM[24980] + MEM[27330];
assign MEM[30871] = MEM[24982] + MEM[25892];
assign MEM[30872] = MEM[24983] + MEM[28967];
assign MEM[30873] = MEM[24985] + MEM[25859];
assign MEM[30874] = MEM[24987] + MEM[28454];
assign MEM[30875] = MEM[24988] + MEM[26586];
assign MEM[30876] = MEM[24990] + MEM[25422];
assign MEM[30877] = MEM[24992] + MEM[25339];
assign MEM[30878] = MEM[24993] + MEM[27585];
assign MEM[30879] = MEM[24994] + MEM[26803];
assign MEM[30880] = MEM[24995] + MEM[27102];
assign MEM[30881] = MEM[24998] + MEM[26554];
assign MEM[30882] = MEM[25000] + MEM[25429];
assign MEM[30883] = MEM[25001] + MEM[26023];
assign MEM[30884] = MEM[25002] + MEM[26473];
assign MEM[30885] = MEM[25005] + MEM[25252];
assign MEM[30886] = MEM[25006] + MEM[26456];
assign MEM[30887] = MEM[25008] + MEM[26340];
assign MEM[30888] = MEM[25010] + MEM[28457];
assign MEM[30889] = MEM[25011] + MEM[27581];
assign MEM[30890] = MEM[25013] + MEM[25288];
assign MEM[30891] = MEM[25017] + MEM[25295];
assign MEM[30892] = MEM[25019] + MEM[26446];
assign MEM[30893] = MEM[25020] + MEM[26667];
assign MEM[30894] = MEM[25021] + MEM[25926];
assign MEM[30895] = MEM[25022] + MEM[28110];
assign MEM[30896] = MEM[25025] + MEM[26893];
assign MEM[30897] = MEM[25026] + MEM[25445];
assign MEM[30898] = MEM[25027] + MEM[25548];
assign MEM[30899] = MEM[25029] + MEM[25516];
assign MEM[30900] = MEM[25030] + MEM[25469];
assign MEM[30901] = MEM[25036] + MEM[26538];
assign MEM[30902] = MEM[25040] + MEM[29334];
assign MEM[30903] = MEM[25045] + MEM[25541];
assign MEM[30904] = MEM[25046] + MEM[26393];
assign MEM[30905] = MEM[25047] + MEM[26530];
assign MEM[30906] = MEM[25049] + MEM[25759];
assign MEM[30907] = MEM[25050] + MEM[27995];
assign MEM[30908] = MEM[25051] + MEM[28072];
assign MEM[30909] = MEM[25052] + MEM[25717];
assign MEM[30910] = MEM[25056] + MEM[27290];
assign MEM[30911] = MEM[25058] + MEM[26302];
assign MEM[30912] = MEM[25059] + MEM[26153];
assign MEM[30913] = MEM[25062] + MEM[26821];
assign MEM[30914] = MEM[25063] + MEM[27138];
assign MEM[30915] = MEM[25064] + MEM[28419];
assign MEM[30916] = MEM[25065] + MEM[25460];
assign MEM[30917] = MEM[25066] + MEM[29987];
assign MEM[30918] = MEM[25067] + MEM[26765];
assign MEM[30919] = MEM[25068] + MEM[26060];
assign MEM[30920] = MEM[25070] + MEM[28225];
assign MEM[30921] = MEM[25072] + MEM[25416];
assign MEM[30922] = MEM[25074] + MEM[25658];
assign MEM[30923] = MEM[25075] + MEM[28991];
assign MEM[30924] = MEM[25077] + MEM[27056];
assign MEM[30925] = MEM[25078] + MEM[28268];
assign MEM[30926] = MEM[25079] + MEM[26733];
assign MEM[30927] = MEM[25080] + MEM[26933];
assign MEM[30928] = MEM[25081] + MEM[29164];
assign MEM[30929] = MEM[25082] + MEM[28036];
assign MEM[30930] = MEM[25083] + MEM[25827];
assign MEM[30931] = MEM[25084] + MEM[28296];
assign MEM[30932] = MEM[25085] + MEM[30318];
assign MEM[30933] = MEM[25088] + MEM[27668];
assign MEM[30934] = MEM[25090] + MEM[27254];
assign MEM[30935] = MEM[25091] + MEM[27665];
assign MEM[30936] = MEM[25092] + MEM[26118];
assign MEM[30937] = MEM[25095] + MEM[27353];
assign MEM[30938] = MEM[25096] + MEM[26024];
assign MEM[30939] = MEM[25097] + MEM[27136];
assign MEM[30940] = MEM[25098] + MEM[26615];
assign MEM[30941] = MEM[25103] + MEM[28990];
assign MEM[30942] = MEM[25104] + MEM[29477];
assign MEM[30943] = MEM[25105] + MEM[25821];
assign MEM[30944] = MEM[25106] + MEM[25508];
assign MEM[30945] = MEM[25107] + MEM[26144];
assign MEM[30946] = MEM[25109] + MEM[26564];
assign MEM[30947] = MEM[25110] + MEM[27270];
assign MEM[30948] = MEM[25111] + MEM[25404];
assign MEM[30949] = MEM[25112] + MEM[26218];
assign MEM[30950] = MEM[25113] + MEM[27486];
assign MEM[30951] = MEM[25114] + MEM[28638];
assign MEM[30952] = MEM[25115] + MEM[29116];
assign MEM[30953] = MEM[25116] + MEM[25355];
assign MEM[30954] = MEM[25117] + MEM[26231];
assign MEM[30955] = MEM[25120] + MEM[26363];
assign MEM[30956] = MEM[25123] + MEM[26661];
assign MEM[30957] = MEM[25127] + MEM[26030];
assign MEM[30958] = MEM[25128] + MEM[25770];
assign MEM[30959] = MEM[25131] + MEM[27403];
assign MEM[30960] = MEM[25133] + MEM[25787];
assign MEM[30961] = MEM[25134] + MEM[27457];
assign MEM[30962] = MEM[25135] + MEM[27480];
assign MEM[30963] = MEM[25137] + MEM[27603];
assign MEM[30964] = MEM[25139] + MEM[27546];
assign MEM[30965] = MEM[25140] + MEM[27708];
assign MEM[30966] = MEM[25142] + MEM[27365];
assign MEM[30967] = MEM[25144] + MEM[26748];
assign MEM[30968] = MEM[25145] + MEM[25836];
assign MEM[30969] = MEM[25146] + MEM[27350];
assign MEM[30970] = MEM[25147] + MEM[25553];
assign MEM[30971] = MEM[25148] + MEM[27049];
assign MEM[30972] = MEM[25151] + MEM[25702];
assign MEM[30973] = MEM[25153] + MEM[25663];
assign MEM[30974] = MEM[25154] + MEM[26464];
assign MEM[30975] = MEM[25156] + MEM[25767];
assign MEM[30976] = MEM[25157] + MEM[27856];
assign MEM[30977] = MEM[25158] + MEM[25897];
assign MEM[30978] = MEM[25159] + MEM[26544];
assign MEM[30979] = MEM[25160] + MEM[25741];
assign MEM[30980] = MEM[25162] + MEM[27649];
assign MEM[30981] = MEM[25164] + MEM[27347];
assign MEM[30982] = MEM[25168] + MEM[26427];
assign MEM[30983] = MEM[25171] + MEM[26912];
assign MEM[30984] = MEM[25172] + MEM[26345];
assign MEM[30985] = MEM[25179] + MEM[29523];
assign MEM[30986] = MEM[25181] + MEM[26262];
assign MEM[30987] = MEM[25183] + MEM[25858];
assign MEM[30988] = MEM[25184] + MEM[27694];
assign MEM[30989] = MEM[25185] + MEM[25559];
assign MEM[30990] = MEM[25196] + MEM[25468];
assign MEM[30991] = MEM[25203] + MEM[26398];
assign MEM[30992] = MEM[25204] + MEM[25626];
assign MEM[30993] = MEM[25205] + MEM[27293];
assign MEM[30994] = MEM[25206] + MEM[26405];
assign MEM[30995] = MEM[25210] + MEM[26179];
assign MEM[30996] = MEM[25211] + MEM[26003];
assign MEM[30997] = MEM[25212] + MEM[27821];
assign MEM[30998] = MEM[25213] + MEM[28720];
assign MEM[30999] = MEM[25214] + MEM[27130];
assign MEM[31000] = MEM[25215] + MEM[25782];
assign MEM[31001] = MEM[25216] + MEM[26284];
assign MEM[31002] = MEM[25217] + MEM[26208];
assign MEM[31003] = MEM[25218] + MEM[27523];
assign MEM[31004] = MEM[25219] + MEM[26533];
assign MEM[31005] = MEM[25220] + MEM[25981];
assign MEM[31006] = MEM[25221] + MEM[26970];
assign MEM[31007] = MEM[25223] + MEM[25577];
assign MEM[31008] = MEM[25224] + MEM[25848];
assign MEM[31009] = MEM[25226] + MEM[26368];
assign MEM[31010] = MEM[25229] + MEM[25539];
assign MEM[31011] = MEM[25231] + MEM[30181];
assign MEM[31012] = MEM[25232] + MEM[26238];
assign MEM[31013] = MEM[25235] + MEM[26362];
assign MEM[31014] = MEM[25236] + MEM[28381];
assign MEM[31015] = MEM[25240] + MEM[27464];
assign MEM[31016] = MEM[25242] + MEM[28764];
assign MEM[31017] = MEM[25243] + MEM[27439];
assign MEM[31018] = MEM[25244] + MEM[28848];
assign MEM[31019] = MEM[25245] + MEM[26745];
assign MEM[31020] = MEM[25246] + MEM[27135];
assign MEM[31021] = MEM[25247] + MEM[26289];
assign MEM[31022] = MEM[25249] + MEM[26267];
assign MEM[31023] = MEM[25250] + MEM[27430];
assign MEM[31024] = MEM[25254] + MEM[26829];
assign MEM[31025] = MEM[25255] + MEM[27466];
assign MEM[31026] = MEM[25256] + MEM[25990];
assign MEM[31027] = MEM[25260] + MEM[26756];
assign MEM[31028] = MEM[25261] + MEM[27530];
assign MEM[31029] = MEM[25262] + MEM[28934];
assign MEM[31030] = MEM[25264] + MEM[25829];
assign MEM[31031] = MEM[25265] + MEM[26654];
assign MEM[31032] = MEM[25267] + MEM[27604];
assign MEM[31033] = MEM[25268] + MEM[26806];
assign MEM[31034] = MEM[25269] + MEM[25845];
assign MEM[31035] = MEM[25272] + MEM[28870];
assign MEM[31036] = MEM[25273] + MEM[26122];
assign MEM[31037] = MEM[25280] + MEM[27499];
assign MEM[31038] = MEM[25282] + MEM[26512];
assign MEM[31039] = MEM[25286] + MEM[28025];
assign MEM[31040] = MEM[25289] + MEM[28952];
assign MEM[31041] = MEM[25292] + MEM[27702];
assign MEM[31042] = MEM[25293] + MEM[27767];
assign MEM[31043] = MEM[25294] + MEM[26753];
assign MEM[31044] = MEM[25296] + MEM[29448];
assign MEM[31045] = MEM[25297] + MEM[26965];
assign MEM[31046] = MEM[25300] + MEM[28485];
assign MEM[31047] = MEM[25301] + MEM[27781];
assign MEM[31048] = MEM[25303] + MEM[27378];
assign MEM[31049] = MEM[25305] + MEM[27268];
assign MEM[31050] = MEM[25306] + MEM[26501];
assign MEM[31051] = MEM[25307] + MEM[25680];
assign MEM[31052] = MEM[25308] + MEM[26998];
assign MEM[31053] = MEM[25309] + MEM[26820];
assign MEM[31054] = MEM[25312] + MEM[25969];
assign MEM[31055] = MEM[25317] + MEM[25977];
assign MEM[31056] = MEM[25320] + MEM[29464];
assign MEM[31057] = MEM[25321] + MEM[25527];
assign MEM[31058] = MEM[25323] + MEM[27375];
assign MEM[31059] = MEM[25324] + MEM[29065];
assign MEM[31060] = MEM[25325] + MEM[29191];
assign MEM[31061] = MEM[25328] + MEM[27876];
assign MEM[31062] = MEM[25329] + MEM[27391];
assign MEM[31063] = MEM[25330] + MEM[27281];
assign MEM[31064] = MEM[25332] + MEM[25784];
assign MEM[31065] = MEM[25333] + MEM[26656];
assign MEM[31066] = MEM[25335] + MEM[26851];
assign MEM[31067] = MEM[25338] + MEM[27490];
assign MEM[31068] = MEM[25340] + MEM[26173];
assign MEM[31069] = MEM[25341] + MEM[25960];
assign MEM[31070] = MEM[25342] + MEM[25885];
assign MEM[31071] = MEM[25343] + MEM[29101];
assign MEM[31072] = MEM[25344] + MEM[26444];
assign MEM[31073] = MEM[25347] + MEM[28335];
assign MEM[31074] = MEM[25348] + MEM[27575];
assign MEM[31075] = MEM[25349] + MEM[27025];
assign MEM[31076] = MEM[25350] + MEM[28620];
assign MEM[31077] = MEM[25351] + MEM[26306];
assign MEM[31078] = MEM[25354] + MEM[28862];
assign MEM[31079] = MEM[25356] + MEM[25943];
assign MEM[31080] = MEM[25357] + MEM[25822];
assign MEM[31081] = MEM[25361] + MEM[26434];
assign MEM[31082] = MEM[25363] + MEM[27363];
assign MEM[31083] = MEM[25365] + MEM[29182];
assign MEM[31084] = MEM[25369] + MEM[26276];
assign MEM[31085] = MEM[25371] + MEM[25800];
assign MEM[31086] = MEM[25372] + MEM[27653];
assign MEM[31087] = MEM[25378] + MEM[25853];
assign MEM[31088] = MEM[25381] + MEM[26072];
assign MEM[31089] = MEM[25384] + MEM[28334];
assign MEM[31090] = MEM[25385] + MEM[26790];
assign MEM[31091] = MEM[25386] + MEM[26561];
assign MEM[31092] = MEM[25387] + MEM[26054];
assign MEM[31093] = MEM[25388] + MEM[26519];
assign MEM[31094] = MEM[25390] + MEM[27073];
assign MEM[31095] = MEM[25391] + MEM[25919];
assign MEM[31096] = MEM[25392] + MEM[27046];
assign MEM[31097] = MEM[25395] + MEM[27300];
assign MEM[31098] = MEM[25396] + MEM[28704];
assign MEM[31099] = MEM[25397] + MEM[28872];
assign MEM[31100] = MEM[25401] + MEM[25463];
assign MEM[31101] = MEM[25403] + MEM[28194];
assign MEM[31102] = MEM[25409] + MEM[26190];
assign MEM[31103] = MEM[25411] + MEM[26201];
assign MEM[31104] = MEM[25412] + MEM[26511];
assign MEM[31105] = MEM[25414] + MEM[26089];
assign MEM[31106] = MEM[25415] + MEM[29072];
assign MEM[31107] = MEM[25423] + MEM[26280];
assign MEM[31108] = MEM[25424] + MEM[26084];
assign MEM[31109] = MEM[25426] + MEM[27001];
assign MEM[31110] = MEM[25427] + MEM[28780];
assign MEM[31111] = MEM[25431] + MEM[28015];
assign MEM[31112] = MEM[25434] + MEM[26429];
assign MEM[31113] = MEM[25435] + MEM[26959];
assign MEM[31114] = MEM[25436] + MEM[25781];
assign MEM[31115] = MEM[25439] + MEM[25844];
assign MEM[31116] = MEM[25441] + MEM[26426];
assign MEM[31117] = MEM[25442] + MEM[26035];
assign MEM[31118] = MEM[25443] + MEM[25584];
assign MEM[31119] = MEM[25446] + MEM[26936];
assign MEM[31120] = MEM[25447] + MEM[29736];
assign MEM[31121] = MEM[25448] + MEM[27654];
assign MEM[31122] = MEM[25449] + MEM[25872];
assign MEM[31123] = MEM[25451] + MEM[25792];
assign MEM[31124] = MEM[25453] + MEM[27823];
assign MEM[31125] = MEM[25454] + MEM[26540];
assign MEM[31126] = MEM[25455] + MEM[27390];
assign MEM[31127] = MEM[25456] + MEM[28427];
assign MEM[31128] = MEM[25462] + MEM[26705];
assign MEM[31129] = MEM[25465] + MEM[30572];
assign MEM[31130] = MEM[25466] + MEM[26780];
assign MEM[31131] = MEM[25467] + MEM[26675];
assign MEM[31132] = MEM[25471] + MEM[28829];
assign MEM[31133] = MEM[25473] + MEM[27178];
assign MEM[31134] = MEM[25475] + MEM[27977];
assign MEM[31135] = MEM[25477] + MEM[27848];
assign MEM[31136] = MEM[25479] + MEM[26197];
assign MEM[31137] = MEM[25480] + MEM[26019];
assign MEM[31138] = MEM[25482] + MEM[29231];
assign MEM[31139] = MEM[25484] + MEM[28912];
assign MEM[31140] = MEM[25485] + MEM[27081];
assign MEM[31141] = MEM[25487] + MEM[26877];
assign MEM[31142] = MEM[25491] + MEM[26835];
assign MEM[31143] = MEM[25494] + MEM[26639];
assign MEM[31144] = MEM[25497] + MEM[29022];
assign MEM[31145] = MEM[25498] + MEM[26277];
assign MEM[31146] = MEM[25499] + MEM[27412];
assign MEM[31147] = MEM[25503] + MEM[25903];
assign MEM[31148] = MEM[25504] + MEM[27671];
assign MEM[31149] = MEM[25505] + MEM[27574];
assign MEM[31150] = MEM[25507] + MEM[26660];
assign MEM[31151] = MEM[25510] + MEM[30577];
assign MEM[31152] = MEM[25511] + MEM[25837];
assign MEM[31153] = MEM[25512] + MEM[29655];
assign MEM[31154] = MEM[25518] + MEM[28784];
assign MEM[31155] = MEM[25520] + MEM[27045];
assign MEM[31156] = MEM[25521] + MEM[25931];
assign MEM[31157] = MEM[25522] + MEM[27108];
assign MEM[31158] = MEM[25524] + MEM[26809];
assign MEM[31159] = MEM[25526] + MEM[26016];
assign MEM[31160] = MEM[25529] + MEM[26138];
assign MEM[31161] = MEM[25530] + MEM[27887];
assign MEM[31162] = MEM[25531] + MEM[28534];
assign MEM[31163] = MEM[25532] + MEM[26924];
assign MEM[31164] = MEM[25534] + MEM[27939];
assign MEM[31165] = MEM[25536] + MEM[27444];
assign MEM[31166] = MEM[25537] + MEM[27518];
assign MEM[31167] = MEM[25538] + MEM[25779];
assign MEM[31168] = MEM[25545] + MEM[28675];
assign MEM[31169] = MEM[25546] + MEM[28440];
assign MEM[31170] = MEM[25547] + MEM[26357];
assign MEM[31171] = MEM[25549] + MEM[26160];
assign MEM[31172] = MEM[25551] + MEM[28265];
assign MEM[31173] = MEM[25552] + MEM[29972];
assign MEM[31174] = MEM[25555] + MEM[27256];
assign MEM[31175] = MEM[25556] + MEM[29216];
assign MEM[31176] = MEM[25560] + MEM[28512];
assign MEM[31177] = MEM[25561] + MEM[27798];
assign MEM[31178] = MEM[25562] + MEM[27311];
assign MEM[31179] = MEM[25564] + MEM[25841];
assign MEM[31180] = MEM[25569] + MEM[26847];
assign MEM[31181] = MEM[25570] + MEM[27866];
assign MEM[31182] = MEM[25571] + MEM[28342];
assign MEM[31183] = MEM[25572] + MEM[30253];
assign MEM[31184] = MEM[25574] + MEM[26369];
assign MEM[31185] = MEM[25575] + MEM[26290];
assign MEM[31186] = MEM[25576] + MEM[25762];
assign MEM[31187] = MEM[25582] + MEM[27777];
assign MEM[31188] = MEM[25585] + MEM[26500];
assign MEM[31189] = MEM[25586] + MEM[28597];
assign MEM[31190] = MEM[25591] + MEM[27213];
assign MEM[31191] = MEM[25595] + MEM[26071];
assign MEM[31192] = MEM[25600] + MEM[26958];
assign MEM[31193] = MEM[25601] + MEM[26477];
assign MEM[31194] = MEM[25603] + MEM[27062];
assign MEM[31195] = MEM[25604] + MEM[26623];
assign MEM[31196] = MEM[25605] + MEM[25920];
assign MEM[31197] = MEM[25608] + MEM[28114];
assign MEM[31198] = MEM[25609] + MEM[26771];
assign MEM[31199] = MEM[25610] + MEM[26181];
assign MEM[31200] = MEM[25611] + MEM[26247];
assign MEM[31201] = MEM[25612] + MEM[25693];
assign MEM[31202] = MEM[25613] + MEM[27113];
assign MEM[31203] = MEM[25614] + MEM[30371];
assign MEM[31204] = MEM[25615] + MEM[26742];
assign MEM[31205] = MEM[25616] + MEM[27435];
assign MEM[31206] = MEM[25617] + MEM[27631];
assign MEM[31207] = MEM[25618] + MEM[27018];
assign MEM[31208] = MEM[25620] + MEM[26739];
assign MEM[31209] = MEM[25621] + MEM[27074];
assign MEM[31210] = MEM[25623] + MEM[26018];
assign MEM[31211] = MEM[25625] + MEM[26752];
assign MEM[31212] = MEM[25627] + MEM[29257];
assign MEM[31213] = MEM[25629] + MEM[27139];
assign MEM[31214] = MEM[25630] + MEM[27874];
assign MEM[31215] = MEM[25631] + MEM[27042];
assign MEM[31216] = MEM[25632] + MEM[27790];
assign MEM[31217] = MEM[25634] + MEM[26228];
assign MEM[31218] = MEM[25636] + MEM[28085];
assign MEM[31219] = MEM[25637] + MEM[27070];
assign MEM[31220] = MEM[25638] + MEM[26269];
assign MEM[31221] = MEM[25639] + MEM[28365];
assign MEM[31222] = MEM[25640] + MEM[26713];
assign MEM[31223] = MEM[25642] + MEM[29251];
assign MEM[31224] = MEM[25643] + MEM[26432];
assign MEM[31225] = MEM[25645] + MEM[25958];
assign MEM[31226] = MEM[25646] + MEM[25899];
assign MEM[31227] = MEM[25647] + MEM[26674];
assign MEM[31228] = MEM[25649] + MEM[27497];
assign MEM[31229] = MEM[25650] + MEM[25839];
assign MEM[31230] = MEM[25652] + MEM[27584];
assign MEM[31231] = MEM[25653] + MEM[27519];
assign MEM[31232] = MEM[25657] + MEM[26333];
assign MEM[31233] = MEM[25659] + MEM[27267];
assign MEM[31234] = MEM[25660] + MEM[25838];
assign MEM[31235] = MEM[25661] + MEM[29275];
assign MEM[31236] = MEM[25664] + MEM[28231];
assign MEM[31237] = MEM[25667] + MEM[26824];
assign MEM[31238] = MEM[25668] + MEM[29033];
assign MEM[31239] = MEM[25669] + MEM[25995];
assign MEM[31240] = MEM[25670] + MEM[26439];
assign MEM[31241] = MEM[25674] + MEM[26701];
assign MEM[31242] = MEM[25675] + MEM[28148];
assign MEM[31243] = MEM[25677] + MEM[29194];
assign MEM[31244] = MEM[25678] + MEM[27638];
assign MEM[31245] = MEM[25681] + MEM[30448];
assign MEM[31246] = MEM[25686] + MEM[29946];
assign MEM[31247] = MEM[25688] + MEM[27847];
assign MEM[31248] = MEM[25689] + MEM[30060];
assign MEM[31249] = MEM[25690] + MEM[29400];
assign MEM[31250] = MEM[25697] + MEM[26596];
assign MEM[31251] = MEM[25700] + MEM[27472];
assign MEM[31252] = MEM[25701] + MEM[26645];
assign MEM[31253] = MEM[25703] + MEM[26609];
assign MEM[31254] = MEM[25704] + MEM[26365];
assign MEM[31255] = MEM[25705] + MEM[26182];
assign MEM[31256] = MEM[25710] + MEM[27532];
assign MEM[31257] = MEM[25712] + MEM[26746];
assign MEM[31258] = MEM[25713] + MEM[26343];
assign MEM[31259] = MEM[25714] + MEM[26879];
assign MEM[31260] = MEM[25716] + MEM[26021];
assign MEM[31261] = MEM[25721] + MEM[27822];
assign MEM[31262] = MEM[25724] + MEM[27468];
assign MEM[31263] = MEM[25725] + MEM[27454];
assign MEM[31264] = MEM[25731] + MEM[27623];
assign MEM[31265] = MEM[25733] + MEM[29359];
assign MEM[31266] = MEM[25735] + MEM[26599];
assign MEM[31267] = MEM[25736] + MEM[27085];
assign MEM[31268] = MEM[25737] + MEM[26066];
assign MEM[31269] = MEM[25738] + MEM[30007];
assign MEM[31270] = MEM[25740] + MEM[29577];
assign MEM[31271] = MEM[25742] + MEM[26625];
assign MEM[31272] = MEM[25748] + MEM[26469];
assign MEM[31273] = MEM[25749] + MEM[28379];
assign MEM[31274] = MEM[25750] + MEM[26584];
assign MEM[31275] = MEM[25752] + MEM[26676];
assign MEM[31276] = MEM[25753] + MEM[29945];
assign MEM[31277] = MEM[25754] + MEM[29195];
assign MEM[31278] = MEM[25756] + MEM[28593];
assign MEM[31279] = MEM[25758] + MEM[28513];
assign MEM[31280] = MEM[25760] + MEM[27151];
assign MEM[31281] = MEM[25763] + MEM[26136];
assign MEM[31282] = MEM[25764] + MEM[27105];
assign MEM[31283] = MEM[25765] + MEM[30020];
assign MEM[31284] = MEM[25766] + MEM[27075];
assign MEM[31285] = MEM[25768] + MEM[28144];
assign MEM[31286] = MEM[25769] + MEM[26960];
assign MEM[31287] = MEM[25777] + MEM[28366];
assign MEM[31288] = MEM[25778] + MEM[27280];
assign MEM[31289] = MEM[25780] + MEM[27424];
assign MEM[31290] = MEM[25783] + MEM[26568];
assign MEM[31291] = MEM[25790] + MEM[29046];
assign MEM[31292] = MEM[25791] + MEM[25986];
assign MEM[31293] = MEM[25793] + MEM[27679];
assign MEM[31294] = MEM[25795] + MEM[26757];
assign MEM[31295] = MEM[25796] + MEM[27912];
assign MEM[31296] = MEM[25797] + MEM[26137];
assign MEM[31297] = MEM[25798] + MEM[28851];
assign MEM[31298] = MEM[25799] + MEM[26589];
assign MEM[31299] = MEM[25802] + MEM[30450];
assign MEM[31300] = MEM[25805] + MEM[27832];
assign MEM[31301] = MEM[25809] + MEM[26031];
assign MEM[31302] = MEM[25811] + MEM[26559];
assign MEM[31303] = MEM[25813] + MEM[27793];
assign MEM[31304] = MEM[25819] + MEM[26775];
assign MEM[31305] = MEM[25823] + MEM[26260];
assign MEM[31306] = MEM[25824] + MEM[26447];
assign MEM[31307] = MEM[25826] + MEM[27014];
assign MEM[31308] = MEM[25828] + MEM[28587];
assign MEM[31309] = MEM[25830] + MEM[29514];
assign MEM[31310] = MEM[25831] + MEM[27415];
assign MEM[31311] = MEM[25832] + MEM[29816];
assign MEM[31312] = MEM[25834] + MEM[26462];
assign MEM[31313] = MEM[25835] + MEM[27937];
assign MEM[31314] = MEM[25840] + MEM[26150];
assign MEM[31315] = MEM[25846] + MEM[28473];
assign MEM[31316] = MEM[25847] + MEM[27508];
assign MEM[31317] = MEM[25852] + MEM[27630];
assign MEM[31318] = MEM[25857] + MEM[27251];
assign MEM[31319] = MEM[25860] + MEM[27644];
assign MEM[31320] = MEM[25864] + MEM[27381];
assign MEM[31321] = MEM[25866] + MEM[28568];
assign MEM[31322] = MEM[25867] + MEM[28140];
assign MEM[31323] = MEM[25868] + MEM[27580];
assign MEM[31324] = MEM[25869] + MEM[30839];
assign MEM[31325] = MEM[25874] + MEM[29110];
assign MEM[31326] = MEM[25876] + MEM[27641];
assign MEM[31327] = MEM[25879] + MEM[29554];
assign MEM[31328] = MEM[25880] + MEM[26579];
assign MEM[31329] = MEM[25884] + MEM[27147];
assign MEM[31330] = MEM[25887] + MEM[27206];
assign MEM[31331] = MEM[25890] + MEM[26935];
assign MEM[31332] = MEM[25894] + MEM[26773];
assign MEM[31333] = MEM[25900] + MEM[28488];
assign MEM[31334] = MEM[25902] + MEM[26092];
assign MEM[31335] = MEM[25904] + MEM[26454];
assign MEM[31336] = MEM[25905] + MEM[27481];
assign MEM[31337] = MEM[25906] + MEM[27167];
assign MEM[31338] = MEM[25907] + MEM[26984];
assign MEM[31339] = MEM[25908] + MEM[27691];
assign MEM[31340] = MEM[25913] + MEM[28936];
assign MEM[31341] = MEM[25915] + MEM[27315];
assign MEM[31342] = MEM[25918] + MEM[28254];
assign MEM[31343] = MEM[25922] + MEM[29529];
assign MEM[31344] = MEM[25924] + MEM[30139];
assign MEM[31345] = MEM[25927] + MEM[29967];
assign MEM[31346] = MEM[25929] + MEM[26367];
assign MEM[31347] = MEM[25933] + MEM[26743];
assign MEM[31348] = MEM[25934] + MEM[30891];
assign MEM[31349] = MEM[25935] + MEM[29380];
assign MEM[31350] = MEM[25937] + MEM[26401];
assign MEM[31351] = MEM[25938] + MEM[29279];
assign MEM[31352] = MEM[25940] + MEM[27080];
assign MEM[31353] = MEM[25941] + MEM[26418];
assign MEM[31354] = MEM[25945] + MEM[26975];
assign MEM[31355] = MEM[25946] + MEM[29151];
assign MEM[31356] = MEM[25949] + MEM[27112];
assign MEM[31357] = MEM[25951] + MEM[29530];
assign MEM[31358] = MEM[25952] + MEM[27714];
assign MEM[31359] = MEM[25954] + MEM[30830];
assign MEM[31360] = MEM[25955] + MEM[27259];
assign MEM[31361] = MEM[25956] + MEM[26891];
assign MEM[31362] = MEM[25962] + MEM[29867];
assign MEM[31363] = MEM[25963] + MEM[29607];
assign MEM[31364] = MEM[25964] + MEM[27098];
assign MEM[31365] = MEM[25965] + MEM[27013];
assign MEM[31366] = MEM[25966] + MEM[27819];
assign MEM[31367] = MEM[25971] + MEM[27160];
assign MEM[31368] = MEM[25972] + MEM[27512];
assign MEM[31369] = MEM[25973] + MEM[26973];
assign MEM[31370] = MEM[25974] + MEM[27205];
assign MEM[31371] = MEM[25975] + MEM[26969];
assign MEM[31372] = MEM[25978] + MEM[27438];
assign MEM[31373] = MEM[25979] + MEM[28075];
assign MEM[31374] = MEM[25982] + MEM[27667];
assign MEM[31375] = MEM[25983] + MEM[26823];
assign MEM[31376] = MEM[25985] + MEM[28565];
assign MEM[31377] = MEM[25987] + MEM[27501];
assign MEM[31378] = MEM[25989] + MEM[27416];
assign MEM[31379] = MEM[25991] + MEM[28792];
assign MEM[31380] = MEM[25993] + MEM[26241];
assign MEM[31381] = MEM[25994] + MEM[26976];
assign MEM[31382] = MEM[25997] + MEM[27560];
assign MEM[31383] = MEM[25998] + MEM[27063];
assign MEM[31384] = MEM[26000] + MEM[26814];
assign MEM[31385] = MEM[26002] + MEM[26598];
assign MEM[31386] = MEM[26004] + MEM[27340];
assign MEM[31387] = MEM[26005] + MEM[26608];
assign MEM[31388] = MEM[26014] + MEM[27297];
assign MEM[31389] = MEM[26026] + MEM[28774];
assign MEM[31390] = MEM[26028] + MEM[27037];
assign MEM[31391] = MEM[26032] + MEM[27789];
assign MEM[31392] = MEM[26034] + MEM[27323];
assign MEM[31393] = MEM[26036] + MEM[27170];
assign MEM[31394] = MEM[26039] + MEM[30082];
assign MEM[31395] = MEM[26043] + MEM[27882];
assign MEM[31396] = MEM[26044] + MEM[27405];
assign MEM[31397] = MEM[26046] + MEM[27142];
assign MEM[31398] = MEM[26047] + MEM[27706];
assign MEM[31399] = MEM[26049] + MEM[26652];
assign MEM[31400] = MEM[26050] + MEM[29036];
assign MEM[31401] = MEM[26051] + MEM[27283];
assign MEM[31402] = MEM[26052] + MEM[27536];
assign MEM[31403] = MEM[26053] + MEM[30493];
assign MEM[31404] = MEM[26055] + MEM[28929];
assign MEM[31405] = MEM[26056] + MEM[28486];
assign MEM[31406] = MEM[26057] + MEM[29541];
assign MEM[31407] = MEM[26059] + MEM[29954];
assign MEM[31408] = MEM[26062] + MEM[26232];
assign MEM[31409] = MEM[26063] + MEM[29265];
assign MEM[31410] = MEM[26064] + MEM[27860];
assign MEM[31411] = MEM[26065] + MEM[27463];
assign MEM[31412] = MEM[26069] + MEM[29354];
assign MEM[31413] = MEM[26070] + MEM[30506];
assign MEM[31414] = MEM[26079] + MEM[27614];
assign MEM[31415] = MEM[26080] + MEM[28372];
assign MEM[31416] = MEM[26082] + MEM[26679];
assign MEM[31417] = MEM[26083] + MEM[30668];
assign MEM[31418] = MEM[26086] + MEM[29677];
assign MEM[31419] = MEM[26088] + MEM[27133];
assign MEM[31420] = MEM[26090] + MEM[30781];
assign MEM[31421] = MEM[26093] + MEM[29537];
assign MEM[31422] = MEM[26094] + MEM[28553];
assign MEM[31423] = MEM[26096] + MEM[26940];
assign MEM[31424] = MEM[26097] + MEM[26419];
assign MEM[31425] = MEM[26098] + MEM[27646];
assign MEM[31426] = MEM[26100] + MEM[28892];
assign MEM[31427] = MEM[26101] + MEM[27816];
assign MEM[31428] = MEM[26102] + MEM[26952];
assign MEM[31429] = MEM[26103] + MEM[27551];
assign MEM[31430] = MEM[26104] + MEM[27906];
assign MEM[31431] = MEM[26106] + MEM[28107];
assign MEM[31432] = MEM[26107] + MEM[27752];
assign MEM[31433] = MEM[26109] + MEM[26431];
assign MEM[31434] = MEM[26111] + MEM[28221];
assign MEM[31435] = MEM[26114] + MEM[28969];
assign MEM[31436] = MEM[26115] + MEM[26458];
assign MEM[31437] = MEM[26117] + MEM[29909];
assign MEM[31438] = MEM[26125] + MEM[28924];
assign MEM[31439] = MEM[26126] + MEM[27813];
assign MEM[31440] = MEM[26128] + MEM[27524];
assign MEM[31441] = MEM[26134] + MEM[27652];
assign MEM[31442] = MEM[26135] + MEM[29578];
assign MEM[31443] = MEM[26141] + MEM[27935];
assign MEM[31444] = MEM[26148] + MEM[28814];
assign MEM[31445] = MEM[26151] + MEM[27513];
assign MEM[31446] = MEM[26152] + MEM[26977];
assign MEM[31447] = MEM[26154] + MEM[27968];
assign MEM[31448] = MEM[26155] + MEM[27885];
assign MEM[31449] = MEM[26158] + MEM[28034];
assign MEM[31450] = MEM[26159] + MEM[27199];
assign MEM[31451] = MEM[26162] + MEM[27202];
assign MEM[31452] = MEM[26163] + MEM[28722];
assign MEM[31453] = MEM[26166] + MEM[28484];
assign MEM[31454] = MEM[26169] + MEM[29528];
assign MEM[31455] = MEM[26172] + MEM[28298];
assign MEM[31456] = MEM[26174] + MEM[29835];
assign MEM[31457] = MEM[26177] + MEM[30700];
assign MEM[31458] = MEM[26178] + MEM[28127];
assign MEM[31459] = MEM[26180] + MEM[27941];
assign MEM[31460] = MEM[26187] + MEM[31234];
assign MEM[31461] = MEM[26188] + MEM[27540];
assign MEM[31462] = MEM[26189] + MEM[27355];
assign MEM[31463] = MEM[26193] + MEM[27775];
assign MEM[31464] = MEM[26196] + MEM[28124];
assign MEM[31465] = MEM[26198] + MEM[27778];
assign MEM[31466] = MEM[26199] + MEM[28639];
assign MEM[31467] = MEM[26200] + MEM[26768];
assign MEM[31468] = MEM[26202] + MEM[29758];
assign MEM[31469] = MEM[26204] + MEM[27181];
assign MEM[31470] = MEM[26209] + MEM[27277];
assign MEM[31471] = MEM[26210] + MEM[29060];
assign MEM[31472] = MEM[26211] + MEM[27159];
assign MEM[31473] = MEM[26212] + MEM[27312];
assign MEM[31474] = MEM[26213] + MEM[27655];
assign MEM[31475] = MEM[26214] + MEM[27372];
assign MEM[31476] = MEM[26216] + MEM[28377];
assign MEM[31477] = MEM[26217] + MEM[29517];
assign MEM[31478] = MEM[26220] + MEM[27361];
assign MEM[31479] = MEM[26221] + MEM[27748];
assign MEM[31480] = MEM[26222] + MEM[26414];
assign MEM[31481] = MEM[26224] + MEM[27388];
assign MEM[31482] = MEM[26226] + MEM[27701];
assign MEM[31483] = MEM[26227] + MEM[30369];
assign MEM[31484] = MEM[26233] + MEM[29080];
assign MEM[31485] = MEM[26234] + MEM[28161];
assign MEM[31486] = MEM[26235] + MEM[27052];
assign MEM[31487] = MEM[26236] + MEM[28008];
assign MEM[31488] = MEM[26237] + MEM[27682];
assign MEM[31489] = MEM[26244] + MEM[27971];
assign MEM[31490] = MEM[26245] + MEM[27455];
assign MEM[31491] = MEM[26248] + MEM[27275];
assign MEM[31492] = MEM[26251] + MEM[28834];
assign MEM[31493] = MEM[26252] + MEM[27828];
assign MEM[31494] = MEM[26254] + MEM[29208];
assign MEM[31495] = MEM[26257] + MEM[28420];
assign MEM[31496] = MEM[26258] + MEM[27418];
assign MEM[31497] = MEM[26264] + MEM[30330];
assign MEM[31498] = MEM[26270] + MEM[27707];
assign MEM[31499] = MEM[26272] + MEM[30164];
assign MEM[31500] = MEM[26273] + MEM[26602];
assign MEM[31501] = MEM[26275] + MEM[27012];
assign MEM[31502] = MEM[26279] + MEM[28563];
assign MEM[31503] = MEM[26282] + MEM[26982];
assign MEM[31504] = MEM[26283] + MEM[28643];
assign MEM[31505] = MEM[26287] + MEM[27924];
assign MEM[31506] = MEM[26292] + MEM[29035];
assign MEM[31507] = MEM[26294] + MEM[27504];
assign MEM[31508] = MEM[26295] + MEM[28061];
assign MEM[31509] = MEM[26296] + MEM[26856];
assign MEM[31510] = MEM[26297] + MEM[28517];
assign MEM[31511] = MEM[26298] + MEM[29198];
assign MEM[31512] = MEM[26299] + MEM[27333];
assign MEM[31513] = MEM[26300] + MEM[26987];
assign MEM[31514] = MEM[26301] + MEM[29652];
assign MEM[31515] = MEM[26303] + MEM[28353];
assign MEM[31516] = MEM[26304] + MEM[29053];
assign MEM[31517] = MEM[26305] + MEM[29152];
assign MEM[31518] = MEM[26307] + MEM[27802];
assign MEM[31519] = MEM[26308] + MEM[26992];
assign MEM[31520] = MEM[26309] + MEM[27367];
assign MEM[31521] = MEM[26314] + MEM[26631];
assign MEM[31522] = MEM[26315] + MEM[26673];
assign MEM[31523] = MEM[26319] + MEM[28132];
assign MEM[31524] = MEM[26322] + MEM[27285];
assign MEM[31525] = MEM[26323] + MEM[29202];
assign MEM[31526] = MEM[26325] + MEM[26878];
assign MEM[31527] = MEM[26326] + MEM[29627];
assign MEM[31528] = MEM[26327] + MEM[27071];
assign MEM[31529] = MEM[26330] + MEM[29190];
assign MEM[31530] = MEM[26332] + MEM[29187];
assign MEM[31531] = MEM[26336] + MEM[29701];
assign MEM[31532] = MEM[26338] + MEM[27855];
assign MEM[31533] = MEM[26339] + MEM[27053];
assign MEM[31534] = MEM[26341] + MEM[28180];
assign MEM[31535] = MEM[26344] + MEM[27296];
assign MEM[31536] = MEM[26346] + MEM[29849];
assign MEM[31537] = MEM[26347] + MEM[27730];
assign MEM[31538] = MEM[26348] + MEM[27534];
assign MEM[31539] = MEM[26349] + MEM[26665];
assign MEM[31540] = MEM[26353] + MEM[27358];
assign MEM[31541] = MEM[26356] + MEM[29425];
assign MEM[31542] = MEM[26359] + MEM[27252];
assign MEM[31543] = MEM[26360] + MEM[27258];
assign MEM[31544] = MEM[26364] + MEM[28113];
assign MEM[31545] = MEM[26374] + MEM[30593];
assign MEM[31546] = MEM[26377] + MEM[28320];
assign MEM[31547] = MEM[26380] + MEM[28893];
assign MEM[31548] = MEM[26384] + MEM[27461];
assign MEM[31549] = MEM[26385] + MEM[27165];
assign MEM[31550] = MEM[26386] + MEM[27209];
assign MEM[31551] = MEM[26387] + MEM[29865];
assign MEM[31552] = MEM[26389] + MEM[27780];
assign MEM[31553] = MEM[26390] + MEM[27015];
assign MEM[31554] = MEM[26395] + MEM[27493];
assign MEM[31555] = MEM[26396] + MEM[28617];
assign MEM[31556] = MEM[26399] + MEM[27492];
assign MEM[31557] = MEM[26400] + MEM[28539];
assign MEM[31558] = MEM[26402] + MEM[26710];
assign MEM[31559] = MEM[26408] + MEM[27891];
assign MEM[31560] = MEM[26409] + MEM[28679];
assign MEM[31561] = MEM[26411] + MEM[26749];
assign MEM[31562] = MEM[26412] + MEM[30527];
assign MEM[31563] = MEM[26413] + MEM[29952];
assign MEM[31564] = MEM[26416] + MEM[27635];
assign MEM[31565] = MEM[26420] + MEM[29158];
assign MEM[31566] = MEM[26421] + MEM[27904];
assign MEM[31567] = MEM[26422] + MEM[27549];
assign MEM[31568] = MEM[26423] + MEM[29707];
assign MEM[31569] = MEM[26424] + MEM[26827];
assign MEM[31570] = MEM[26425] + MEM[28903];
assign MEM[31571] = MEM[26428] + MEM[28219];
assign MEM[31572] = MEM[26430] + MEM[30691];
assign MEM[31573] = MEM[26433] + MEM[27969];
assign MEM[31574] = MEM[26437] + MEM[28826];
assign MEM[31575] = MEM[26440] + MEM[27208];
assign MEM[31576] = MEM[26445] + MEM[28515];
assign MEM[31577] = MEM[26450] + MEM[26776];
assign MEM[31578] = MEM[26451] + MEM[27915];
assign MEM[31579] = MEM[26453] + MEM[28843];
assign MEM[31580] = MEM[26457] + MEM[27506];
assign MEM[31581] = MEM[26463] + MEM[27253];
assign MEM[31582] = MEM[26466] + MEM[26968];
assign MEM[31583] = MEM[26470] + MEM[28044];
assign MEM[31584] = MEM[26472] + MEM[27769];
assign MEM[31585] = MEM[26474] + MEM[26647];
assign MEM[31586] = MEM[26475] + MEM[30949];
assign MEM[31587] = MEM[26476] + MEM[27782];
assign MEM[31588] = MEM[26479] + MEM[26557];
assign MEM[31589] = MEM[26482] + MEM[27035];
assign MEM[31590] = MEM[26487] + MEM[30057];
assign MEM[31591] = MEM[26490] + MEM[27121];
assign MEM[31592] = MEM[26492] + MEM[26777];
assign MEM[31593] = MEM[26493] + MEM[30672];
assign MEM[31594] = MEM[26496] + MEM[29715];
assign MEM[31595] = MEM[26498] + MEM[27899];
assign MEM[31596] = MEM[26502] + MEM[28845];
assign MEM[31597] = MEM[26503] + MEM[28619];
assign MEM[31598] = MEM[26506] + MEM[27449];
assign MEM[31599] = MEM[26507] + MEM[30234];
assign MEM[31600] = MEM[26508] + MEM[30362];
assign MEM[31601] = MEM[26513] + MEM[29281];
assign MEM[31602] = MEM[26514] + MEM[27568];
assign MEM[31603] = MEM[26515] + MEM[27236];
assign MEM[31604] = MEM[26517] + MEM[27970];
assign MEM[31605] = MEM[26518] + MEM[26761];
assign MEM[31606] = MEM[26520] + MEM[26655];
assign MEM[31607] = MEM[26521] + MEM[30132];
assign MEM[31608] = MEM[26522] + MEM[28039];
assign MEM[31609] = MEM[26524] + MEM[27043];
assign MEM[31610] = MEM[26527] + MEM[28658];
assign MEM[31611] = MEM[26528] + MEM[27966];
assign MEM[31612] = MEM[26529] + MEM[27547];
assign MEM[31613] = MEM[26531] + MEM[29067];
assign MEM[31614] = MEM[26534] + MEM[28198];
assign MEM[31615] = MEM[26536] + MEM[28269];
assign MEM[31616] = MEM[26537] + MEM[26868];
assign MEM[31617] = MEM[26539] + MEM[30957];
assign MEM[31618] = MEM[26542] + MEM[26772];
assign MEM[31619] = MEM[26543] + MEM[29884];
assign MEM[31620] = MEM[26546] + MEM[30512];
assign MEM[31621] = MEM[26548] + MEM[27997];
assign MEM[31622] = MEM[26550] + MEM[28183];
assign MEM[31623] = MEM[26551] + MEM[27441];
assign MEM[31624] = MEM[26556] + MEM[27910];
assign MEM[31625] = MEM[26558] + MEM[27685];
assign MEM[31626] = MEM[26560] + MEM[28744];
assign MEM[31627] = MEM[26562] + MEM[30605];
assign MEM[31628] = MEM[26565] + MEM[27677];
assign MEM[31629] = MEM[26567] + MEM[27166];
assign MEM[31630] = MEM[26569] + MEM[28552];
assign MEM[31631] = MEM[26571] + MEM[28333];
assign MEM[31632] = MEM[26573] + MEM[27599];
assign MEM[31633] = MEM[26574] + MEM[29001];
assign MEM[31634] = MEM[26576] + MEM[27800];
assign MEM[31635] = MEM[26580] + MEM[27739];
assign MEM[31636] = MEM[26581] + MEM[27397];
assign MEM[31637] = MEM[26582] + MEM[28166];
assign MEM[31638] = MEM[26583] + MEM[27693];
assign MEM[31639] = MEM[26585] + MEM[27784];
assign MEM[31640] = MEM[26592] + MEM[27741];
assign MEM[31641] = MEM[26594] + MEM[29520];
assign MEM[31642] = MEM[26595] + MEM[27619];
assign MEM[31643] = MEM[26600] + MEM[28806];
assign MEM[31644] = MEM[26601] + MEM[30412];
assign MEM[31645] = MEM[26603] + MEM[29658];
assign MEM[31646] = MEM[26605] + MEM[28582];
assign MEM[31647] = MEM[26606] + MEM[29282];
assign MEM[31648] = MEM[26613] + MEM[28385];
assign MEM[31649] = MEM[26614] + MEM[27284];
assign MEM[31650] = MEM[26616] + MEM[30312];
assign MEM[31651] = MEM[26618] + MEM[30152];
assign MEM[31652] = MEM[26620] + MEM[28948];
assign MEM[31653] = MEM[26622] + MEM[27522];
assign MEM[31654] = MEM[26627] + MEM[27187];
assign MEM[31655] = MEM[26628] + MEM[28038];
assign MEM[31656] = MEM[26629] + MEM[27842];
assign MEM[31657] = MEM[26630] + MEM[27527];
assign MEM[31658] = MEM[26632] + MEM[28270];
assign MEM[31659] = MEM[26633] + MEM[27692];
assign MEM[31660] = MEM[26634] + MEM[27651];
assign MEM[31661] = MEM[26635] + MEM[27379];
assign MEM[31662] = MEM[26636] + MEM[28088];
assign MEM[31663] = MEM[26637] + MEM[29654];
assign MEM[31664] = MEM[26638] + MEM[26895];
assign MEM[31665] = MEM[26640] + MEM[27398];
assign MEM[31666] = MEM[26641] + MEM[31145];
assign MEM[31667] = MEM[26642] + MEM[29792];
assign MEM[31668] = MEM[26643] + MEM[28153];
assign MEM[31669] = MEM[26653] + MEM[27624];
assign MEM[31670] = MEM[26657] + MEM[29196];
assign MEM[31671] = MEM[26658] + MEM[28491];
assign MEM[31672] = MEM[26663] + MEM[29699];
assign MEM[31673] = MEM[26666] + MEM[30693];
assign MEM[31674] = MEM[26668] + MEM[27109];
assign MEM[31675] = MEM[26669] + MEM[28817];
assign MEM[31676] = MEM[26670] + MEM[27395];
assign MEM[31677] = MEM[26671] + MEM[27786];
assign MEM[31678] = MEM[26672] + MEM[28271];
assign MEM[31679] = MEM[26680] + MEM[29525];
assign MEM[31680] = MEM[26681] + MEM[29019];
assign MEM[31681] = MEM[26684] + MEM[27020];
assign MEM[31682] = MEM[26685] + MEM[28559];
assign MEM[31683] = MEM[26687] + MEM[30484];
assign MEM[31684] = MEM[26690] + MEM[28984];
assign MEM[31685] = MEM[26691] + MEM[30843];
assign MEM[31686] = MEM[26692] + MEM[28625];
assign MEM[31687] = MEM[26693] + MEM[28621];
assign MEM[31688] = MEM[26694] + MEM[27409];
assign MEM[31689] = MEM[26695] + MEM[28395];
assign MEM[31690] = MEM[26696] + MEM[28229];
assign MEM[31691] = MEM[26697] + MEM[28048];
assign MEM[31692] = MEM[26698] + MEM[30513];
assign MEM[31693] = MEM[26699] + MEM[27510];
assign MEM[31694] = MEM[26700] + MEM[27943];
assign MEM[31695] = MEM[26703] + MEM[28476];
assign MEM[31696] = MEM[26708] + MEM[27172];
assign MEM[31697] = MEM[26709] + MEM[27389];
assign MEM[31698] = MEM[26714] + MEM[27385];
assign MEM[31699] = MEM[26715] + MEM[28536];
assign MEM[31700] = MEM[26717] + MEM[27859];
assign MEM[31701] = MEM[26719] + MEM[29798];
assign MEM[31702] = MEM[26721] + MEM[27716];
assign MEM[31703] = MEM[26723] + MEM[28078];
assign MEM[31704] = MEM[26724] + MEM[30452];
assign MEM[31705] = MEM[26726] + MEM[27442];
assign MEM[31706] = MEM[26728] + MEM[31050];
assign MEM[31707] = MEM[26731] + MEM[28329];
assign MEM[31708] = MEM[26732] + MEM[28650];
assign MEM[31709] = MEM[26734] + MEM[27201];
assign MEM[31710] = MEM[26735] + MEM[27950];
assign MEM[31711] = MEM[26736] + MEM[28428];
assign MEM[31712] = MEM[26737] + MEM[29340];
assign MEM[31713] = MEM[26738] + MEM[27414];
assign MEM[31714] = MEM[26741] + MEM[30345];
assign MEM[31715] = MEM[26747] + MEM[27198];
assign MEM[31716] = MEM[26754] + MEM[28055];
assign MEM[31717] = MEM[26755] + MEM[28607];
assign MEM[31718] = MEM[26763] + MEM[28277];
assign MEM[31719] = MEM[26764] + MEM[27994];
assign MEM[31720] = MEM[26766] + MEM[28331];
assign MEM[31721] = MEM[26770] + MEM[30106];
assign MEM[31722] = MEM[26774] + MEM[30215];
assign MEM[31723] = MEM[26779] + MEM[29968];
assign MEM[31724] = MEM[26781] + MEM[27705];
assign MEM[31725] = MEM[26783] + MEM[29268];
assign MEM[31726] = MEM[26786] + MEM[28742];
assign MEM[31727] = MEM[26791] + MEM[28453];
assign MEM[31728] = MEM[26793] + MEM[28600];
assign MEM[31729] = MEM[26794] + MEM[28528];
assign MEM[31730] = MEM[26795] + MEM[27550];
assign MEM[31731] = MEM[26796] + MEM[30143];
assign MEM[31732] = MEM[26797] + MEM[30198];
assign MEM[31733] = MEM[26799] + MEM[28226];
assign MEM[31734] = MEM[26800] + MEM[27925];
assign MEM[31735] = MEM[26810] + MEM[29088];
assign MEM[31736] = MEM[26813] + MEM[29511];
assign MEM[31737] = MEM[26816] + MEM[28199];
assign MEM[31738] = MEM[26817] + MEM[29238];
assign MEM[31739] = MEM[26819] + MEM[29572];
assign MEM[31740] = MEM[26822] + MEM[29727];
assign MEM[31741] = MEM[26825] + MEM[28024];
assign MEM[31742] = MEM[26826] + MEM[29481];
assign MEM[31743] = MEM[26828] + MEM[28137];
assign MEM[31744] = MEM[26830] + MEM[27945];
assign MEM[31745] = MEM[26832] + MEM[28416];
assign MEM[31746] = MEM[26834] + MEM[29171];
assign MEM[31747] = MEM[26837] + MEM[30069];
assign MEM[31748] = MEM[26838] + MEM[28546];
assign MEM[31749] = MEM[26839] + MEM[30171];
assign MEM[31750] = MEM[26840] + MEM[28781];
assign MEM[31751] = MEM[26842] + MEM[29333];
assign MEM[31752] = MEM[26843] + MEM[28500];
assign MEM[31753] = MEM[26844] + MEM[29555];
assign MEM[31754] = MEM[26845] + MEM[28407];
assign MEM[31755] = MEM[26846] + MEM[27586];
assign MEM[31756] = MEM[26848] + MEM[29762];
assign MEM[31757] = MEM[26849] + MEM[28212];
assign MEM[31758] = MEM[26850] + MEM[30677];
assign MEM[31759] = MEM[26853] + MEM[27661];
assign MEM[31760] = MEM[26855] + MEM[29714];
assign MEM[31761] = MEM[26858] + MEM[30800];
assign MEM[31762] = MEM[26859] + MEM[29133];
assign MEM[31763] = MEM[26861] + MEM[28927];
assign MEM[31764] = MEM[26862] + MEM[29249];
assign MEM[31765] = MEM[26863] + MEM[29348];
assign MEM[31766] = MEM[26864] + MEM[27681];
assign MEM[31767] = MEM[26865] + MEM[27091];
assign MEM[31768] = MEM[26866] + MEM[28431];
assign MEM[31769] = MEM[26867] + MEM[27342];
assign MEM[31770] = MEM[26869] + MEM[29959];
assign MEM[31771] = MEM[26870] + MEM[27124];
assign MEM[31772] = MEM[26871] + MEM[28672];
assign MEM[31773] = MEM[26872] + MEM[27036];
assign MEM[31774] = MEM[26873] + MEM[30533];
assign MEM[31775] = MEM[26875] + MEM[29587];
assign MEM[31776] = MEM[26876] + MEM[27229];
assign MEM[31777] = MEM[26882] + MEM[27875];
assign MEM[31778] = MEM[26883] + MEM[28202];
assign MEM[31779] = MEM[26885] + MEM[27470];
assign MEM[31780] = MEM[26886] + MEM[29252];
assign MEM[31781] = MEM[26887] + MEM[28721];
assign MEM[31782] = MEM[26889] + MEM[29543];
assign MEM[31783] = MEM[26892] + MEM[27920];
assign MEM[31784] = MEM[26894] + MEM[29905];
assign MEM[31785] = MEM[26898] + MEM[27469];
assign MEM[31786] = MEM[26899] + MEM[29512];
assign MEM[31787] = MEM[26904] + MEM[30938];
assign MEM[31788] = MEM[26906] + MEM[28423];
assign MEM[31789] = MEM[26907] + MEM[30737];
assign MEM[31790] = MEM[26909] + MEM[27690];
assign MEM[31791] = MEM[26910] + MEM[29621];
assign MEM[31792] = MEM[26911] + MEM[27615];
assign MEM[31793] = MEM[26914] + MEM[29592];
assign MEM[31794] = MEM[26916] + MEM[30333];
assign MEM[31795] = MEM[26917] + MEM[27407];
assign MEM[31796] = MEM[26920] + MEM[31199];
assign MEM[31797] = MEM[26921] + MEM[29698];
assign MEM[31798] = MEM[26923] + MEM[30204];
assign MEM[31799] = MEM[26925] + MEM[28414];
assign MEM[31800] = MEM[26926] + MEM[27660];
assign MEM[31801] = MEM[26928] + MEM[29866];
assign MEM[31802] = MEM[26931] + MEM[29199];
assign MEM[31803] = MEM[26932] + MEM[27984];
assign MEM[31804] = MEM[26937] + MEM[27485];
assign MEM[31805] = MEM[26938] + MEM[29516];
assign MEM[31806] = MEM[26939] + MEM[27726];
assign MEM[31807] = MEM[26942] + MEM[30372];
assign MEM[31808] = MEM[26943] + MEM[28677];
assign MEM[31809] = MEM[26944] + MEM[28013];
assign MEM[31810] = MEM[26945] + MEM[28752];
assign MEM[31811] = MEM[26946] + MEM[30392];
assign MEM[31812] = MEM[26947] + MEM[30504];
assign MEM[31813] = MEM[26948] + MEM[28820];
assign MEM[31814] = MEM[26949] + MEM[29802];
assign MEM[31815] = MEM[26950] + MEM[28810];
assign MEM[31816] = MEM[26951] + MEM[30380];
assign MEM[31817] = MEM[26953] + MEM[28404];
assign MEM[31818] = MEM[26954] + MEM[28010];
assign MEM[31819] = MEM[26956] + MEM[28685];
assign MEM[31820] = MEM[26957] + MEM[30425];
assign MEM[31821] = MEM[26961] + MEM[27176];
assign MEM[31822] = MEM[26963] + MEM[30034];
assign MEM[31823] = MEM[26966] + MEM[27642];
assign MEM[31824] = MEM[26967] + MEM[28637];
assign MEM[31825] = MEM[26971] + MEM[28095];
assign MEM[31826] = MEM[26972] + MEM[30156];
assign MEM[31827] = MEM[26974] + MEM[29790];
assign MEM[31828] = MEM[26981] + MEM[28782];
assign MEM[31829] = MEM[26985] + MEM[27905];
assign MEM[31830] = MEM[26986] + MEM[29407];
assign MEM[31831] = MEM[26988] + MEM[30000];
assign MEM[31832] = MEM[26989] + MEM[29634];
assign MEM[31833] = MEM[26990] + MEM[28317];
assign MEM[31834] = MEM[26991] + MEM[29963];
assign MEM[31835] = MEM[26993] + MEM[29665];
assign MEM[31836] = MEM[26994] + MEM[28710];
assign MEM[31837] = MEM[26995] + MEM[30765];
assign MEM[31838] = MEM[26996] + MEM[28895];
assign MEM[31839] = MEM[26997] + MEM[27608];
assign MEM[31840] = MEM[27000] + MEM[27543];
assign MEM[31841] = MEM[27002] + MEM[30537];
assign MEM[31842] = MEM[27003] + MEM[27672];
assign MEM[31843] = MEM[27004] + MEM[29519];
assign MEM[31844] = MEM[27006] + MEM[28719];
assign MEM[31845] = MEM[27008] + MEM[28983];
assign MEM[31846] = MEM[27009] + MEM[27721];
assign MEM[31847] = MEM[27010] + MEM[27533];
assign MEM[31848] = MEM[27011] + MEM[29601];
assign MEM[31849] = MEM[27017] + MEM[28158];
assign MEM[31850] = MEM[27021] + MEM[27735];
assign MEM[31851] = MEM[27023] + MEM[29419];
assign MEM[31852] = MEM[27026] + MEM[29939];
assign MEM[31853] = MEM[27027] + MEM[27964];
assign MEM[31854] = MEM[27029] + MEM[27503];
assign MEM[31855] = MEM[27030] + MEM[28472];
assign MEM[31856] = MEM[27032] + MEM[27380];
assign MEM[31857] = MEM[27033] + MEM[28471];
assign MEM[31858] = MEM[27039] + MEM[28739];
assign MEM[31859] = MEM[27040] + MEM[29211];
assign MEM[31860] = MEM[27041] + MEM[27827];
assign MEM[31861] = MEM[27044] + MEM[30612];
assign MEM[31862] = MEM[27048] + MEM[29585];
assign MEM[31863] = MEM[27050] + MEM[28045];
assign MEM[31864] = MEM[27051] + MEM[30273];
assign MEM[31865] = MEM[27057] + MEM[28557];
assign MEM[31866] = MEM[27059] + MEM[30460];
assign MEM[31867] = MEM[27061] + MEM[29825];
assign MEM[31868] = MEM[27064] + MEM[28383];
assign MEM[31869] = MEM[27065] + MEM[27565];
assign MEM[31870] = MEM[27067] + MEM[28059];
assign MEM[31871] = MEM[27068] + MEM[27433];
assign MEM[31872] = MEM[27077] + MEM[27230];
assign MEM[31873] = MEM[27079] + MEM[27628];
assign MEM[31874] = MEM[27082] + MEM[28728];
assign MEM[31875] = MEM[27084] + MEM[28394];
assign MEM[31876] = MEM[27086] + MEM[30240];
assign MEM[31877] = MEM[27088] + MEM[27940];
assign MEM[31878] = MEM[27089] + MEM[27369];
assign MEM[31879] = MEM[27092] + MEM[28009];
assign MEM[31880] = MEM[27094] + MEM[28411];
assign MEM[31881] = MEM[27095] + MEM[29289];
assign MEM[31882] = MEM[27096] + MEM[28823];
assign MEM[31883] = MEM[27097] + MEM[29619];
assign MEM[31884] = MEM[27099] + MEM[27933];
assign MEM[31885] = MEM[27101] + MEM[30269];
assign MEM[31886] = MEM[27103] + MEM[28855];
assign MEM[31887] = MEM[27104] + MEM[29375];
assign MEM[31888] = MEM[27106] + MEM[27772];
assign MEM[31889] = MEM[27107] + MEM[30747];
assign MEM[31890] = MEM[27111] + MEM[30280];
assign MEM[31891] = MEM[27114] + MEM[27958];
assign MEM[31892] = MEM[27115] + MEM[27411];
assign MEM[31893] = MEM[27116] + MEM[29157];
assign MEM[31894] = MEM[27117] + MEM[27851];
assign MEM[31895] = MEM[27119] + MEM[29461];
assign MEM[31896] = MEM[27120] + MEM[30072];
assign MEM[31897] = MEM[27122] + MEM[29146];
assign MEM[31898] = MEM[27123] + MEM[30219];
assign MEM[31899] = MEM[27128] + MEM[27233];
assign MEM[31900] = MEM[27129] + MEM[29928];
assign MEM[31901] = MEM[27131] + MEM[27476];
assign MEM[31902] = MEM[27132] + MEM[29112];
assign MEM[31903] = MEM[27134] + MEM[27299];
assign MEM[31904] = MEM[27137] + MEM[29524];
assign MEM[31905] = MEM[27140] + MEM[30884];
assign MEM[31906] = MEM[27141] + MEM[30377];
assign MEM[31907] = MEM[27143] + MEM[27548];
assign MEM[31908] = MEM[27144] + MEM[28079];
assign MEM[31909] = MEM[27145] + MEM[30465];
assign MEM[31910] = MEM[27146] + MEM[29623];
assign MEM[31911] = MEM[27153] + MEM[27647];
assign MEM[31912] = MEM[27155] + MEM[27460];
assign MEM[31913] = MEM[27156] + MEM[28313];
assign MEM[31914] = MEM[27157] + MEM[27727];
assign MEM[31915] = MEM[27158] + MEM[28109];
assign MEM[31916] = MEM[27161] + MEM[28797];
assign MEM[31917] = MEM[27162] + MEM[28152];
assign MEM[31918] = MEM[27163] + MEM[28354];
assign MEM[31919] = MEM[27168] + MEM[27765];
assign MEM[31920] = MEM[27169] + MEM[28701];
assign MEM[31921] = MEM[27174] + MEM[28982];
assign MEM[31922] = MEM[27175] + MEM[27858];
assign MEM[31923] = MEM[27177] + MEM[28046];
assign MEM[31924] = MEM[27179] + MEM[27243];
assign MEM[31925] = MEM[27180] + MEM[28598];
assign MEM[31926] = MEM[27182] + MEM[27514];
assign MEM[31927] = MEM[27183] + MEM[30749];
assign MEM[31928] = MEM[27184] + MEM[29062];
assign MEM[31929] = MEM[27186] + MEM[29079];
assign MEM[31930] = MEM[27188] + MEM[29611];
assign MEM[31931] = MEM[27189] + MEM[29129];
assign MEM[31932] = MEM[27190] + MEM[28314];
assign MEM[31933] = MEM[27191] + MEM[28054];
assign MEM[31934] = MEM[27192] + MEM[30287];
assign MEM[31935] = MEM[27194] + MEM[31119];
assign MEM[31936] = MEM[27196] + MEM[28388];
assign MEM[31937] = MEM[27197] + MEM[27505];
assign MEM[31938] = MEM[27203] + MEM[28170];
assign MEM[31939] = MEM[27204] + MEM[30186];
assign MEM[31940] = MEM[27207] + MEM[28712];
assign MEM[31941] = MEM[27210] + MEM[28341];
assign MEM[31942] = MEM[27211] + MEM[30422];
assign MEM[31943] = MEM[27212] + MEM[27478];
assign MEM[31944] = MEM[27215] + MEM[28384];
assign MEM[31945] = MEM[27216] + MEM[27852];
assign MEM[31946] = MEM[27219] + MEM[27462];
assign MEM[31947] = MEM[27220] + MEM[29267];
assign MEM[31948] = MEM[27222] + MEM[28671];
assign MEM[31949] = MEM[27223] + MEM[28303];
assign MEM[31950] = MEM[27224] + MEM[29683];
assign MEM[31951] = MEM[27225] + MEM[30008];
assign MEM[31952] = MEM[27227] + MEM[29304];
assign MEM[31953] = MEM[27228] + MEM[27688];
assign MEM[31954] = MEM[27231] + MEM[28940];
assign MEM[31955] = MEM[27232] + MEM[29343];
assign MEM[31956] = MEM[27234] + MEM[28660];
assign MEM[31957] = MEM[27235] + MEM[28011];
assign MEM[31958] = MEM[27237] + MEM[30265];
assign MEM[31959] = MEM[27238] + MEM[29710];
assign MEM[31960] = MEM[27239] + MEM[28753];
assign MEM[31961] = MEM[27241] + MEM[29105];
assign MEM[31962] = MEM[27242] + MEM[29206];
assign MEM[31963] = MEM[27244] + MEM[27783];
assign MEM[31964] = MEM[27245] + MEM[29459];
assign MEM[31965] = MEM[27246] + MEM[27662];
assign MEM[31966] = MEM[27255] + MEM[29544];
assign MEM[31967] = MEM[27260] + MEM[28935];
assign MEM[31968] = MEM[27264] + MEM[28580];
assign MEM[31969] = MEM[27266] + MEM[28964];
assign MEM[31970] = MEM[27269] + MEM[30226];
assign MEM[31971] = MEM[27271] + MEM[31057];
assign MEM[31972] = MEM[27272] + MEM[31186];
assign MEM[31973] = MEM[27273] + MEM[29155];
assign MEM[31974] = MEM[27274] + MEM[27535];
assign MEM[31975] = MEM[27276] + MEM[29215];
assign MEM[31976] = MEM[27286] + MEM[30449];
assign MEM[31977] = MEM[27288] + MEM[28623];
assign MEM[31978] = MEM[27289] + MEM[28426];
assign MEM[31979] = MEM[27291] + MEM[28437];
assign MEM[31980] = MEM[27292] + MEM[31160];
assign MEM[31981] = MEM[27294] + MEM[27750];
assign MEM[31982] = MEM[27295] + MEM[27903];
assign MEM[31983] = MEM[27301] + MEM[28800];
assign MEM[31984] = MEM[27302] + MEM[29119];
assign MEM[31985] = MEM[27305] + MEM[30588];
assign MEM[31986] = MEM[27306] + MEM[30203];
assign MEM[31987] = MEM[27307] + MEM[27456];
assign MEM[31988] = MEM[27308] + MEM[28415];
assign MEM[31989] = MEM[27309] + MEM[27496];
assign MEM[31990] = MEM[27313] + MEM[27382];
assign MEM[31991] = MEM[27314] + MEM[31184];
assign MEM[31992] = MEM[27316] + MEM[28647];
assign MEM[31993] = MEM[27318] + MEM[28725];
assign MEM[31994] = MEM[27319] + MEM[29663];
assign MEM[31995] = MEM[27321] + MEM[30801];
assign MEM[31996] = MEM[27324] + MEM[27812];
assign MEM[31997] = MEM[27325] + MEM[30356];
assign MEM[31998] = MEM[27326] + MEM[31353];
assign MEM[31999] = MEM[27327] + MEM[29058];
assign MEM[32000] = MEM[27328] + MEM[29285];
assign MEM[32001] = MEM[27331] + MEM[28108];
assign MEM[32002] = MEM[27332] + MEM[28082];
assign MEM[32003] = MEM[27334] + MEM[29974];
assign MEM[32004] = MEM[27336] + MEM[29777];
assign MEM[32005] = MEM[27338] + MEM[28119];
assign MEM[32006] = MEM[27341] + MEM[29754];
assign MEM[32007] = MEM[27343] + MEM[30979];
assign MEM[32008] = MEM[27345] + MEM[29290];
assign MEM[32009] = MEM[27348] + MEM[29311];
assign MEM[32010] = MEM[27354] + MEM[29943];
assign MEM[32011] = MEM[27356] + MEM[28544];
assign MEM[32012] = MEM[27357] + MEM[28363];
assign MEM[32013] = MEM[27359] + MEM[28883];
assign MEM[32014] = MEM[27362] + MEM[30463];
assign MEM[32015] = MEM[27364] + MEM[27963];
assign MEM[32016] = MEM[27366] + MEM[30634];
assign MEM[32017] = MEM[27368] + MEM[28874];
assign MEM[32018] = MEM[27370] + MEM[28121];
assign MEM[32019] = MEM[27373] + MEM[29526];
assign MEM[32020] = MEM[27374] + MEM[28798];
assign MEM[32021] = MEM[27376] + MEM[30217];
assign MEM[32022] = MEM[27377] + MEM[29214];
assign MEM[32023] = MEM[27383] + MEM[28946];
assign MEM[32024] = MEM[27384] + MEM[28974];
assign MEM[32025] = MEM[27387] + MEM[29179];
assign MEM[32026] = MEM[27392] + MEM[28868];
assign MEM[32027] = MEM[27393] + MEM[29402];
assign MEM[32028] = MEM[27399] + MEM[28706];
assign MEM[32029] = MEM[27400] + MEM[29172];
assign MEM[32030] = MEM[27402] + MEM[28130];
assign MEM[32031] = MEM[27404] + MEM[29719];
assign MEM[32032] = MEM[27406] + MEM[28661];
assign MEM[32033] = MEM[27408] + MEM[27927];
assign MEM[32034] = MEM[27413] + MEM[30567];
assign MEM[32035] = MEM[27419] + MEM[27948];
assign MEM[32036] = MEM[27421] + MEM[27583];
assign MEM[32037] = MEM[27423] + MEM[29029];
assign MEM[32038] = MEM[27425] + MEM[28734];
assign MEM[32039] = MEM[27426] + MEM[28456];
assign MEM[32040] = MEM[27427] + MEM[29929];
assign MEM[32041] = MEM[27428] + MEM[27509];
assign MEM[32042] = MEM[27429] + MEM[29466];
assign MEM[32043] = MEM[27431] + MEM[30833];
assign MEM[32044] = MEM[27432] + MEM[27762];
assign MEM[32045] = MEM[27434] + MEM[28378];
assign MEM[32046] = MEM[27436] + MEM[29063];
assign MEM[32047] = MEM[27437] + MEM[27587];
assign MEM[32048] = MEM[27443] + MEM[28645];
assign MEM[32049] = MEM[27445] + MEM[30227];
assign MEM[32050] = MEM[27446] + MEM[28570];
assign MEM[32051] = MEM[27448] + MEM[27829];
assign MEM[32052] = MEM[27450] + MEM[28018];
assign MEM[32053] = MEM[27451] + MEM[29270];
assign MEM[32054] = MEM[27453] + MEM[30112];
assign MEM[32055] = MEM[27458] + MEM[28012];
assign MEM[32056] = MEM[27459] + MEM[27854];
assign MEM[32057] = MEM[27465] + MEM[28663];
assign MEM[32058] = MEM[27467] + MEM[30687];
assign MEM[32059] = MEM[27473] + MEM[31141];
assign MEM[32060] = MEM[27474] + MEM[28432];
assign MEM[32061] = MEM[27475] + MEM[27601];
assign MEM[32062] = MEM[27477] + MEM[30409];
assign MEM[32063] = MEM[27479] + MEM[29642];
assign MEM[32064] = MEM[27482] + MEM[27907];
assign MEM[32065] = MEM[27484] + MEM[28368];
assign MEM[32066] = MEM[27487] + MEM[31022];
assign MEM[32067] = MEM[27488] + MEM[30516];
assign MEM[32068] = MEM[27489] + MEM[28604];
assign MEM[32069] = MEM[27491] + MEM[27787];
assign MEM[32070] = MEM[27494] + MEM[30138];
assign MEM[32071] = MEM[27495] + MEM[29721];
assign MEM[32072] = MEM[27498] + MEM[29839];
assign MEM[32073] = MEM[27500] + MEM[29774];
assign MEM[32074] = MEM[27502] + MEM[28066];
assign MEM[32075] = MEM[27507] + MEM[29876];
assign MEM[32076] = MEM[27511] + MEM[29470];
assign MEM[32077] = MEM[27515] + MEM[29061];
assign MEM[32078] = MEM[27517] + MEM[28696];
assign MEM[32079] = MEM[27520] + MEM[30978];
assign MEM[32080] = MEM[27525] + MEM[30462];
assign MEM[32081] = MEM[27526] + MEM[27754];
assign MEM[32082] = MEM[27528] + MEM[27861];
assign MEM[32083] = MEM[27529] + MEM[27704];
assign MEM[32084] = MEM[27537] + MEM[29596];
assign MEM[32085] = MEM[27538] + MEM[30328];
assign MEM[32086] = MEM[27539] + MEM[28156];
assign MEM[32087] = MEM[27545] + MEM[30930];
assign MEM[32088] = MEM[27552] + MEM[30440];
assign MEM[32089] = MEM[27553] + MEM[30637];
assign MEM[32090] = MEM[27554] + MEM[30073];
assign MEM[32091] = MEM[27555] + MEM[29059];
assign MEM[32092] = MEM[27556] + MEM[30346];
assign MEM[32093] = MEM[27558] + MEM[27799];
assign MEM[32094] = MEM[27561] + MEM[27761];
assign MEM[32095] = MEM[27564] + MEM[28131];
assign MEM[32096] = MEM[27566] + MEM[30819];
assign MEM[32097] = MEM[27567] + MEM[27825];
assign MEM[32098] = MEM[27569] + MEM[27913];
assign MEM[32099] = MEM[27570] + MEM[28689];
assign MEM[32100] = MEM[27571] + MEM[28280];
assign MEM[32101] = MEM[27573] + MEM[30790];
assign MEM[32102] = MEM[27576] + MEM[29484];
assign MEM[32103] = MEM[27577] + MEM[29135];
assign MEM[32104] = MEM[27578] + MEM[29286];
assign MEM[32105] = MEM[27579] + MEM[29978];
assign MEM[32106] = MEM[27589] + MEM[28711];
assign MEM[32107] = MEM[27590] + MEM[29889];
assign MEM[32108] = MEM[27591] + MEM[28462];
assign MEM[32109] = MEM[27592] + MEM[30955];
assign MEM[32110] = MEM[27593] + MEM[28190];
assign MEM[32111] = MEM[27594] + MEM[28337];
assign MEM[32112] = MEM[27595] + MEM[28264];
assign MEM[32113] = MEM[27596] + MEM[28757];
assign MEM[32114] = MEM[27600] + MEM[30602];
assign MEM[32115] = MEM[27602] + MEM[29747];
assign MEM[32116] = MEM[27606] + MEM[30314];
assign MEM[32117] = MEM[27607] + MEM[29542];
assign MEM[32118] = MEM[27609] + MEM[29050];
assign MEM[32119] = MEM[27610] + MEM[27909];
assign MEM[32120] = MEM[27611] + MEM[28105];
assign MEM[32121] = MEM[27612] + MEM[29298];
assign MEM[32122] = MEM[27613] + MEM[28651];
assign MEM[32123] = MEM[27616] + MEM[31393];
assign MEM[32124] = MEM[27617] + MEM[28033];
assign MEM[32125] = MEM[27618] + MEM[28886];
assign MEM[32126] = MEM[27621] + MEM[29391];
assign MEM[32127] = MEM[27622] + MEM[28091];
assign MEM[32128] = MEM[27625] + MEM[28211];
assign MEM[32129] = MEM[27626] + MEM[29264];
assign MEM[32130] = MEM[27627] + MEM[28361];
assign MEM[32131] = MEM[27629] + MEM[30841];
assign MEM[32132] = MEM[27632] + MEM[30053];
assign MEM[32133] = MEM[27633] + MEM[28707];
assign MEM[32134] = MEM[27634] + MEM[27845];
assign MEM[32135] = MEM[27636] + MEM[29538];
assign MEM[32136] = MEM[27637] + MEM[29881];
assign MEM[32137] = MEM[27639] + MEM[28616];
assign MEM[32138] = MEM[27640] + MEM[30650];
assign MEM[32139] = MEM[27643] + MEM[28310];
assign MEM[32140] = MEM[27645] + MEM[31017];
assign MEM[32141] = MEM[27648] + MEM[28525];
assign MEM[32142] = MEM[27657] + MEM[28831];
assign MEM[32143] = MEM[27659] + MEM[28747];
assign MEM[32144] = MEM[27663] + MEM[28740];
assign MEM[32145] = MEM[27666] + MEM[30172];
assign MEM[32146] = MEM[27670] + MEM[30755];
assign MEM[32147] = MEM[27673] + MEM[27804];
assign MEM[32148] = MEM[27674] + MEM[28804];
assign MEM[32149] = MEM[27675] + MEM[30582];
assign MEM[32150] = MEM[27676] + MEM[28057];
assign MEM[32151] = MEM[27678] + MEM[28205];
assign MEM[32152] = MEM[27680] + MEM[29420];
assign MEM[32153] = MEM[27683] + MEM[30308];
assign MEM[32154] = MEM[27684] + MEM[28171];
assign MEM[32155] = MEM[27686] + MEM[27831];
assign MEM[32156] = MEM[27687] + MEM[30080];
assign MEM[32157] = MEM[27689] + MEM[30325];
assign MEM[32158] = MEM[27695] + MEM[31251];
assign MEM[32159] = MEM[27696] + MEM[28586];
assign MEM[32160] = MEM[27697] + MEM[29156];
assign MEM[32161] = MEM[27698] + MEM[28478];
assign MEM[32162] = MEM[27699] + MEM[28896];
assign MEM[32163] = MEM[27700] + MEM[27838];
assign MEM[32164] = MEM[27703] + MEM[29292];
assign MEM[32165] = MEM[27709] + MEM[29457];
assign MEM[32166] = MEM[27710] + MEM[28858];
assign MEM[32167] = MEM[27711] + MEM[29370];
assign MEM[32168] = MEM[27712] + MEM[28255];
assign MEM[32169] = MEM[27713] + MEM[28308];
assign MEM[32170] = MEM[27715] + MEM[28827];
assign MEM[32171] = MEM[27717] + MEM[30329];
assign MEM[32172] = MEM[27718] + MEM[28863];
assign MEM[32173] = MEM[27720] + MEM[28003];
assign MEM[32174] = MEM[27723] + MEM[28899];
assign MEM[32175] = MEM[27724] + MEM[28356];
assign MEM[32176] = MEM[27725] + MEM[31108];
assign MEM[32177] = MEM[27729] + MEM[31210];
assign MEM[32178] = MEM[27731] + MEM[28435];
assign MEM[32179] = MEM[27732] + MEM[27965];
assign MEM[32180] = MEM[27733] + MEM[30803];
assign MEM[32181] = MEM[27734] + MEM[28591];
assign MEM[32182] = MEM[27738] + MEM[30896];
assign MEM[32183] = MEM[27740] + MEM[28309];
assign MEM[32184] = MEM[27742] + MEM[27944];
assign MEM[32185] = MEM[27743] + MEM[31066];
assign MEM[32186] = MEM[27744] + MEM[31033];
assign MEM[32187] = MEM[27745] + MEM[28162];
assign MEM[32188] = MEM[27746] + MEM[31024];
assign MEM[32189] = MEM[27747] + MEM[28588];
assign MEM[32190] = MEM[27749] + MEM[29937];
assign MEM[32191] = MEM[27751] + MEM[29540];
assign MEM[32192] = MEM[27753] + MEM[30569];
assign MEM[32193] = MEM[27755] + MEM[27811];
assign MEM[32194] = MEM[27756] + MEM[28470];
assign MEM[32195] = MEM[27757] + MEM[28956];
assign MEM[32196] = MEM[27758] + MEM[30768];
assign MEM[32197] = MEM[27759] + MEM[31367];
assign MEM[32198] = MEM[27760] + MEM[29923];
assign MEM[32199] = MEM[27763] + MEM[28441];
assign MEM[32200] = MEM[27764] + MEM[31356];
assign MEM[32201] = MEM[27766] + MEM[28509];
assign MEM[32202] = MEM[27768] + MEM[30945];
assign MEM[32203] = MEM[27770] + MEM[28301];
assign MEM[32204] = MEM[27771] + MEM[30868];
assign MEM[32205] = MEM[27773] + MEM[28632];
assign MEM[32206] = MEM[27774] + MEM[28266];
assign MEM[32207] = MEM[27779] + MEM[28708];
assign MEM[32208] = MEM[27785] + MEM[28410];
assign MEM[32209] = MEM[27794] + MEM[28263];
assign MEM[32210] = MEM[27795] + MEM[30247];
assign MEM[32211] = MEM[27796] + MEM[28071];
assign MEM[32212] = MEM[27797] + MEM[30670];
assign MEM[32213] = MEM[27801] + MEM[29506];
assign MEM[32214] = MEM[27803] + MEM[30870];
assign MEM[32215] = MEM[27805] + MEM[29427];
assign MEM[32216] = MEM[27806] + MEM[28325];
assign MEM[32217] = MEM[27807] + MEM[28766];
assign MEM[32218] = MEM[27808] + MEM[28386];
assign MEM[32219] = MEM[27809] + MEM[28538];
assign MEM[32220] = MEM[27810] + MEM[29392];
assign MEM[32221] = MEM[27814] + MEM[30926];
assign MEM[32222] = MEM[27815] + MEM[29643];
assign MEM[32223] = MEM[27817] + MEM[28944];
assign MEM[32224] = MEM[27818] + MEM[28128];
assign MEM[32225] = MEM[27820] + MEM[29097];
assign MEM[32226] = MEM[27824] + MEM[29515];
assign MEM[32227] = MEM[27830] + MEM[28636];
assign MEM[32228] = MEM[27834] + MEM[28216];
assign MEM[32229] = MEM[27835] + MEM[29118];
assign MEM[32230] = MEM[27836] + MEM[28247];
assign MEM[32231] = MEM[27837] + MEM[30108];
assign MEM[32232] = MEM[27839] + MEM[29324];
assign MEM[32233] = MEM[27840] + MEM[28238];
assign MEM[32234] = MEM[27841] + MEM[28041];
assign MEM[32235] = MEM[27843] + MEM[27955];
assign MEM[32236] = MEM[27844] + MEM[30315];
assign MEM[32237] = MEM[27846] + MEM[28052];
assign MEM[32238] = MEM[27849] + MEM[29903];
assign MEM[32239] = MEM[27850] + MEM[28908];
assign MEM[32240] = MEM[27853] + MEM[29647];
assign MEM[32241] = MEM[27857] + MEM[28289];
assign MEM[32242] = MEM[27862] + MEM[30489];
assign MEM[32243] = MEM[27863] + MEM[30962];
assign MEM[32244] = MEM[27864] + MEM[30190];
assign MEM[32245] = MEM[27865] + MEM[28727];
assign MEM[32246] = MEM[27867] + MEM[28434];
assign MEM[32247] = MEM[27868] + MEM[30378];
assign MEM[32248] = MEM[27869] + MEM[31226];
assign MEM[32249] = MEM[27871] + MEM[30148];
assign MEM[32250] = MEM[27872] + MEM[28323];
assign MEM[32251] = MEM[27873] + MEM[31196];
assign MEM[32252] = MEM[27877] + MEM[31094];
assign MEM[32253] = MEM[27878] + MEM[28151];
assign MEM[32254] = MEM[27879] + MEM[30100];
assign MEM[32255] = MEM[27880] + MEM[28291];
assign MEM[32256] = MEM[27883] + MEM[28547];
assign MEM[32257] = MEM[27884] + MEM[28497];
assign MEM[32258] = MEM[27886] + MEM[28535];
assign MEM[32259] = MEM[27888] + MEM[30545];
assign MEM[32260] = MEM[27889] + MEM[28135];
assign MEM[32261] = MEM[27890] + MEM[30578];
assign MEM[32262] = MEM[27892] + MEM[28352];
assign MEM[32263] = MEM[27893] + MEM[28763];
assign MEM[32264] = MEM[27894] + MEM[29123];
assign MEM[32265] = MEM[27895] + MEM[28902];
assign MEM[32266] = MEM[27897] + MEM[28963];
assign MEM[32267] = MEM[27898] + MEM[29416];
assign MEM[32268] = MEM[27900] + MEM[28514];
assign MEM[32269] = MEM[27901] + MEM[29726];
assign MEM[32270] = MEM[27908] + MEM[28228];
assign MEM[32271] = MEM[27911] + MEM[31384];
assign MEM[32272] = MEM[27916] + MEM[29864];
assign MEM[32273] = MEM[27917] + MEM[30393];
assign MEM[32274] = MEM[27918] + MEM[28242];
assign MEM[32275] = MEM[27919] + MEM[28606];
assign MEM[32276] = MEM[27921] + MEM[30405];
assign MEM[32277] = MEM[27922] + MEM[29947];
assign MEM[32278] = MEM[27923] + MEM[29637];
assign MEM[32279] = MEM[27926] + MEM[28795];
assign MEM[32280] = MEM[27928] + MEM[28307];
assign MEM[32281] = MEM[27929] + MEM[29234];
assign MEM[32282] = MEM[27930] + MEM[30004];
assign MEM[32283] = MEM[27931] + MEM[28813];
assign MEM[32284] = MEM[27932] + MEM[29588];
assign MEM[32285] = MEM[27934] + MEM[28001];
assign MEM[32286] = MEM[27938] + MEM[30116];
assign MEM[32287] = MEM[27942] + MEM[28519];
assign MEM[32288] = MEM[27946] + MEM[28771];
assign MEM[32289] = MEM[27947] + MEM[29040];
assign MEM[32290] = MEM[27951] + MEM[29130];
assign MEM[32291] = MEM[27952] + MEM[28890];
assign MEM[32292] = MEM[27953] + MEM[29629];
assign MEM[32293] = MEM[27956] + MEM[30319];
assign MEM[32294] = MEM[27957] + MEM[29349];
assign MEM[32295] = MEM[27959] + MEM[28859];
assign MEM[32296] = MEM[27960] + MEM[28793];
assign MEM[32297] = MEM[27961] + MEM[30821];
assign MEM[32298] = MEM[27962] + MEM[29418];
assign MEM[32299] = MEM[27967] + MEM[28328];
assign MEM[32300] = MEM[27972] + MEM[28168];
assign MEM[32301] = MEM[27973] + MEM[28391];
assign MEM[32302] = MEM[27974] + MEM[29413];
assign MEM[32303] = MEM[27975] + MEM[27998];
assign MEM[32304] = MEM[27976] + MEM[28447];
assign MEM[32305] = MEM[27978] + MEM[30291];
assign MEM[32306] = MEM[27982] + MEM[31003];
assign MEM[32307] = MEM[27983] + MEM[31360];
assign MEM[32308] = MEM[27986] + MEM[28233];
assign MEM[32309] = MEM[27987] + MEM[31028];
assign MEM[32310] = MEM[27989] + MEM[31423];
assign MEM[32311] = MEM[27990] + MEM[30610];
assign MEM[32312] = MEM[27991] + MEM[28175];
assign MEM[32313] = MEM[27993] + MEM[30894];
assign MEM[32314] = MEM[27999] + MEM[29431];
assign MEM[32315] = MEM[28000] + MEM[31539];
assign MEM[32316] = MEM[28002] + MEM[28402];
assign MEM[32317] = MEM[28004] + MEM[30144];
assign MEM[32318] = MEM[28005] + MEM[28550];
assign MEM[32319] = MEM[28006] + MEM[30558];
assign MEM[32320] = MEM[28007] + MEM[28240];
assign MEM[32321] = MEM[28014] + MEM[29789];
assign MEM[32322] = MEM[28016] + MEM[28201];
assign MEM[32323] = MEM[28017] + MEM[29045];
assign MEM[32324] = MEM[28020] + MEM[31581];
assign MEM[32325] = MEM[28022] + MEM[30658];
assign MEM[32326] = MEM[28023] + MEM[29632];
assign MEM[32327] = MEM[28027] + MEM[31364];
assign MEM[32328] = MEM[28029] + MEM[29492];
assign MEM[32329] = MEM[28030] + MEM[28692];
assign MEM[32330] = MEM[28031] + MEM[28717];
assign MEM[32331] = MEM[28032] + MEM[29605];
assign MEM[32332] = MEM[28035] + MEM[28302];
assign MEM[32333] = MEM[28040] + MEM[28421];
assign MEM[32334] = MEM[28042] + MEM[28316];
assign MEM[32335] = MEM[28043] + MEM[31042];
assign MEM[32336] = MEM[28051] + MEM[30353];
assign MEM[32337] = MEM[28053] + MEM[31177];
assign MEM[32338] = MEM[28056] + MEM[29852];
assign MEM[32339] = MEM[28058] + MEM[28567];
assign MEM[32340] = MEM[28060] + MEM[29951];
assign MEM[32341] = MEM[28062] + MEM[29114];
assign MEM[32342] = MEM[28063] + MEM[28665];
assign MEM[32343] = MEM[28064] + MEM[29869];
assign MEM[32344] = MEM[28067] + MEM[28227];
assign MEM[32345] = MEM[28068] + MEM[30370];
assign MEM[32346] = MEM[28069] + MEM[29509];
assign MEM[32347] = MEM[28070] + MEM[30160];
assign MEM[32348] = MEM[28076] + MEM[28173];
assign MEM[32349] = MEM[28080] + MEM[28987];
assign MEM[32350] = MEM[28081] + MEM[30756];
assign MEM[32351] = MEM[28084] + MEM[28724];
assign MEM[32352] = MEM[28086] + MEM[28783];
assign MEM[32353] = MEM[28089] + MEM[30402];
assign MEM[32354] = MEM[28090] + MEM[28479];
assign MEM[32355] = MEM[28092] + MEM[30389];
assign MEM[32356] = MEM[28093] + MEM[28475];
assign MEM[32357] = MEM[28094] + MEM[31304];
assign MEM[32358] = MEM[28096] + MEM[29344];
assign MEM[32359] = MEM[28097] + MEM[29984];
assign MEM[32360] = MEM[28098] + MEM[28844];
assign MEM[32361] = MEM[28099] + MEM[28464];
assign MEM[32362] = MEM[28100] + MEM[28482];
assign MEM[32363] = MEM[28101] + MEM[30381];
assign MEM[32364] = MEM[28103] + MEM[30278];
assign MEM[32365] = MEM[28104] + MEM[28819];
assign MEM[32366] = MEM[28106] + MEM[28501];
assign MEM[32367] = MEM[28111] + MEM[29870];
assign MEM[32368] = MEM[28112] + MEM[29069];
assign MEM[32369] = MEM[28115] + MEM[30736];
assign MEM[32370] = MEM[28117] + MEM[28919];
assign MEM[32371] = MEM[28118] + MEM[31716];
assign MEM[32372] = MEM[28120] + MEM[31642];
assign MEM[32373] = MEM[28122] + MEM[28815];
assign MEM[32374] = MEM[28123] + MEM[29219];
assign MEM[32375] = MEM[28125] + MEM[31187];
assign MEM[32376] = MEM[28126] + MEM[29472];
assign MEM[32377] = MEM[28133] + MEM[28502];
assign MEM[32378] = MEM[28134] + MEM[28345];
assign MEM[32379] = MEM[28138] + MEM[28885];
assign MEM[32380] = MEM[28139] + MEM[28449];
assign MEM[32381] = MEM[28142] + MEM[31638];
assign MEM[32382] = MEM[28143] + MEM[28569];
assign MEM[32383] = MEM[28145] + MEM[31425];
assign MEM[32384] = MEM[28146] + MEM[28718];
assign MEM[32385] = MEM[28147] + MEM[30231];
assign MEM[32386] = MEM[28149] + MEM[30618];
assign MEM[32387] = MEM[28150] + MEM[29934];
assign MEM[32388] = MEM[28155] + MEM[30633];
assign MEM[32389] = MEM[28157] + MEM[28294];
assign MEM[32390] = MEM[28159] + MEM[28733];
assign MEM[32391] = MEM[28163] + MEM[29176];
assign MEM[32392] = MEM[28165] + MEM[30199];
assign MEM[32393] = MEM[28167] + MEM[28408];
assign MEM[32394] = MEM[28169] + MEM[29757];
assign MEM[32395] = MEM[28172] + MEM[31777];
assign MEM[32396] = MEM[28174] + MEM[29042];
assign MEM[32397] = MEM[28176] + MEM[31475];
assign MEM[32398] = MEM[28177] + MEM[32041];
assign MEM[32399] = MEM[28178] + MEM[28397];
assign MEM[32400] = MEM[28179] + MEM[30710];
assign MEM[32401] = MEM[28182] + MEM[28778];
assign MEM[32402] = MEM[28184] + MEM[29183];
assign MEM[32403] = MEM[28185] + MEM[29468];
assign MEM[32404] = MEM[28187] + MEM[29948];
assign MEM[32405] = MEM[28188] + MEM[30078];
assign MEM[32406] = MEM[28192] + MEM[29581];
assign MEM[32407] = MEM[28193] + MEM[28901];
assign MEM[32408] = MEM[28195] + MEM[30151];
assign MEM[32409] = MEM[28196] + MEM[28493];
assign MEM[32410] = MEM[28197] + MEM[28370];
assign MEM[32411] = MEM[28200] + MEM[29617];
assign MEM[32412] = MEM[28203] + MEM[29174];
assign MEM[32413] = MEM[28204] + MEM[29501];
assign MEM[32414] = MEM[28206] + MEM[29443];
assign MEM[32415] = MEM[28207] + MEM[28374];
assign MEM[32416] = MEM[28208] + MEM[29931];
assign MEM[32417] = MEM[28209] + MEM[28678];
assign MEM[32418] = MEM[28210] + MEM[28709];
assign MEM[32419] = MEM[28213] + MEM[31113];
assign MEM[32420] = MEM[28214] + MEM[28686];
assign MEM[32421] = MEM[28215] + MEM[29013];
assign MEM[32422] = MEM[28217] + MEM[29859];
assign MEM[32423] = MEM[28220] + MEM[28847];
assign MEM[32424] = MEM[28222] + MEM[31411];
assign MEM[32425] = MEM[28223] + MEM[31823];
assign MEM[32426] = MEM[28224] + MEM[28581];
assign MEM[32427] = MEM[28232] + MEM[31354];
assign MEM[32428] = MEM[28234] + MEM[29011];
assign MEM[32429] = MEM[28235] + MEM[29661];
assign MEM[32430] = MEM[28236] + MEM[29084];
assign MEM[32431] = MEM[28237] + MEM[28866];
assign MEM[32432] = MEM[28239] + MEM[31263];
assign MEM[32433] = MEM[28241] + MEM[29579];
assign MEM[32434] = MEM[28244] + MEM[30624];
assign MEM[32435] = MEM[28245] + MEM[29393];
assign MEM[32436] = MEM[28246] + MEM[28926];
assign MEM[32437] = MEM[28248] + MEM[29522];
assign MEM[32438] = MEM[28249] + MEM[29955];
assign MEM[32439] = MEM[28250] + MEM[30006];
assign MEM[32440] = MEM[28251] + MEM[29565];
assign MEM[32441] = MEM[28252] + MEM[29606];
assign MEM[32442] = MEM[28253] + MEM[29153];
assign MEM[32443] = MEM[28257] + MEM[31111];
assign MEM[32444] = MEM[28258] + MEM[29310];
assign MEM[32445] = MEM[28259] + MEM[30154];
assign MEM[32446] = MEM[28260] + MEM[31157];
assign MEM[32447] = MEM[28261] + MEM[28433];
assign MEM[32448] = MEM[28262] + MEM[29454];
assign MEM[32449] = MEM[28267] + MEM[28918];
assign MEM[32450] = MEM[28272] + MEM[29969];
assign MEM[32451] = MEM[28273] + MEM[28953];
assign MEM[32452] = MEM[28275] + MEM[29679];
assign MEM[32453] = MEM[28276] + MEM[31715];
assign MEM[32454] = MEM[28278] + MEM[31668];
assign MEM[32455] = MEM[28279] + MEM[29720];
assign MEM[32456] = MEM[28281] + MEM[29192];
assign MEM[32457] = MEM[28282] + MEM[29505];
assign MEM[32458] = MEM[28283] + MEM[31267];
assign MEM[32459] = MEM[28284] + MEM[29007];
assign MEM[32460] = MEM[28285] + MEM[28787];
assign MEM[32461] = MEM[28287] + MEM[30011];
assign MEM[32462] = MEM[28288] + MEM[28424];
assign MEM[32463] = MEM[28290] + MEM[29557];
assign MEM[32464] = MEM[28295] + MEM[30631];
assign MEM[32465] = MEM[28297] + MEM[31259];
assign MEM[32466] = MEM[28299] + MEM[28396];
assign MEM[32467] = MEM[28300] + MEM[29043];
assign MEM[32468] = MEM[28304] + MEM[28799];
assign MEM[32469] = MEM[28305] + MEM[28596];
assign MEM[32470] = MEM[28306] + MEM[31220];
assign MEM[32471] = MEM[28311] + MEM[28676];
assign MEM[32472] = MEM[28312] + MEM[30183];
assign MEM[32473] = MEM[28315] + MEM[30119];
assign MEM[32474] = MEM[28318] + MEM[30548];
assign MEM[32475] = MEM[28319] + MEM[31030];
assign MEM[32476] = MEM[28322] + MEM[29048];
assign MEM[32477] = MEM[28324] + MEM[28654];
assign MEM[32478] = MEM[28327] + MEM[29303];
assign MEM[32479] = MEM[28330] + MEM[30187];
assign MEM[32480] = MEM[28336] + MEM[30161];
assign MEM[32481] = MEM[28338] + MEM[28958];
assign MEM[32482] = MEM[28339] + MEM[28495];
assign MEM[32483] = MEM[28340] + MEM[31149];
assign MEM[32484] = MEM[28343] + MEM[29609];
assign MEM[32485] = MEM[28346] + MEM[30528];
assign MEM[32486] = MEM[28347] + MEM[31290];
assign MEM[32487] = MEM[28348] + MEM[30435];
assign MEM[32488] = MEM[28349] + MEM[31271];
assign MEM[32489] = MEM[28351] + MEM[29186];
assign MEM[32490] = MEM[28355] + MEM[31785];
assign MEM[32491] = MEM[28357] + MEM[29144];
assign MEM[32492] = MEM[28358] + MEM[29269];
assign MEM[32493] = MEM[28359] + MEM[31588];
assign MEM[32494] = MEM[28362] + MEM[31724];
assign MEM[32495] = MEM[28364] + MEM[30763];
assign MEM[32496] = MEM[28367] + MEM[31419];
assign MEM[32497] = MEM[28369] + MEM[30141];
assign MEM[32498] = MEM[28371] + MEM[28670];
assign MEM[32499] = MEM[28376] + MEM[29902];
assign MEM[32500] = MEM[28380] + MEM[31170];
assign MEM[32501] = MEM[28382] + MEM[30754];
assign MEM[32502] = MEM[28387] + MEM[29204];
assign MEM[32503] = MEM[28389] + MEM[29326];
assign MEM[32504] = MEM[28390] + MEM[28659];
assign MEM[32505] = MEM[28393] + MEM[29432];
assign MEM[32506] = MEM[28398] + MEM[30895];
assign MEM[32507] = MEM[28399] + MEM[30867];
assign MEM[32508] = MEM[28400] + MEM[31660];
assign MEM[32509] = MEM[28401] + MEM[29222];
assign MEM[32510] = MEM[28403] + MEM[28429];
assign MEM[32511] = MEM[28405] + MEM[29180];
assign MEM[32512] = MEM[28409] + MEM[28906];
assign MEM[32513] = MEM[28412] + MEM[29589];
assign MEM[32514] = MEM[28413] + MEM[30281];
assign MEM[32515] = MEM[28417] + MEM[30122];
assign MEM[32516] = MEM[28425] + MEM[30214];
assign MEM[32517] = MEM[28430] + MEM[29032];
assign MEM[32518] = MEM[28436] + MEM[29453];
assign MEM[32519] = MEM[28438] + MEM[31681];
assign MEM[32520] = MEM[28445] + MEM[28609];
assign MEM[32521] = MEM[28446] + MEM[29640];
assign MEM[32522] = MEM[28448] + MEM[29189];
assign MEM[32523] = MEM[28450] + MEM[30266];
assign MEM[32524] = MEM[28451] + MEM[31146];
assign MEM[32525] = MEM[28452] + MEM[30505];
assign MEM[32526] = MEM[28455] + MEM[29168];
assign MEM[32527] = MEM[28458] + MEM[30180];
assign MEM[32528] = MEM[28460] + MEM[31609];
assign MEM[32529] = MEM[28461] + MEM[28629];
assign MEM[32530] = MEM[28463] + MEM[28995];
assign MEM[32531] = MEM[28465] + MEM[30804];
assign MEM[32532] = MEM[28467] + MEM[29124];
assign MEM[32533] = MEM[28468] + MEM[30740];
assign MEM[32534] = MEM[28469] + MEM[30288];
assign MEM[32535] = MEM[28474] + MEM[30549];
assign MEM[32536] = MEM[28477] + MEM[30883];
assign MEM[32537] = MEM[28480] + MEM[28888];
assign MEM[32538] = MEM[28481] + MEM[29350];
assign MEM[32539] = MEM[28483] + MEM[29966];
assign MEM[32540] = MEM[28489] + MEM[30350];
assign MEM[32541] = MEM[28490] + MEM[28577];
assign MEM[32542] = MEM[28492] + MEM[32285];
assign MEM[32543] = MEM[28494] + MEM[29412];
assign MEM[32544] = MEM[28496] + MEM[30021];
assign MEM[32545] = MEM[28498] + MEM[30439];
assign MEM[32546] = MEM[28503] + MEM[29496];
assign MEM[32547] = MEM[28505] + MEM[30969];
assign MEM[32548] = MEM[28506] + MEM[30583];
assign MEM[32549] = MEM[28507] + MEM[29729];
assign MEM[32550] = MEM[28508] + MEM[29408];
assign MEM[32551] = MEM[28510] + MEM[29843];
assign MEM[32552] = MEM[28511] + MEM[28558];
assign MEM[32553] = MEM[28516] + MEM[29487];
assign MEM[32554] = MEM[28518] + MEM[30845];
assign MEM[32555] = MEM[28522] + MEM[30245];
assign MEM[32556] = MEM[28526] + MEM[31254];
assign MEM[32557] = MEM[28527] + MEM[30002];
assign MEM[32558] = MEM[28530] + MEM[30968];
assign MEM[32559] = MEM[28531] + MEM[30013];
assign MEM[32560] = MEM[28532] + MEM[28595];
assign MEM[32561] = MEM[28533] + MEM[30262];
assign MEM[32562] = MEM[28537] + MEM[30684];
assign MEM[32563] = MEM[28540] + MEM[29302];
assign MEM[32564] = MEM[28541] + MEM[29965];
assign MEM[32565] = MEM[28542] + MEM[31159];
assign MEM[32566] = MEM[28543] + MEM[30947];
assign MEM[32567] = MEM[28548] + MEM[30097];
assign MEM[32568] = MEM[28549] + MEM[29137];
assign MEM[32569] = MEM[28551] + MEM[30459];
assign MEM[32570] = MEM[28554] + MEM[30596];
assign MEM[32571] = MEM[28556] + MEM[29971];
assign MEM[32572] = MEM[28561] + MEM[31534];
assign MEM[32573] = MEM[28562] + MEM[28773];
assign MEM[32574] = MEM[28564] + MEM[29386];
assign MEM[32575] = MEM[28566] + MEM[30555];
assign MEM[32576] = MEM[28571] + MEM[30935];
assign MEM[32577] = MEM[28572] + MEM[29184];
assign MEM[32578] = MEM[28573] + MEM[29973];
assign MEM[32579] = MEM[28574] + MEM[31391];
assign MEM[32580] = MEM[28575] + MEM[30529];
assign MEM[32581] = MEM[28576] + MEM[29925];
assign MEM[32582] = MEM[28578] + MEM[29141];
assign MEM[32583] = MEM[28579] + MEM[30622];
assign MEM[32584] = MEM[28583] + MEM[29521];
assign MEM[32585] = MEM[28585] + MEM[29761];
assign MEM[32586] = MEM[28589] + MEM[30436];
assign MEM[32587] = MEM[28590] + MEM[28960];
assign MEM[32588] = MEM[28592] + MEM[29668];
assign MEM[32589] = MEM[28594] + MEM[31289];
assign MEM[32590] = MEM[28599] + MEM[28825];
assign MEM[32591] = MEM[28601] + MEM[29560];
assign MEM[32592] = MEM[28602] + MEM[29126];
assign MEM[32593] = MEM[28603] + MEM[30695];
assign MEM[32594] = MEM[28605] + MEM[29574];
assign MEM[32595] = MEM[28608] + MEM[28923];
assign MEM[32596] = MEM[28610] + MEM[30490];
assign MEM[32597] = MEM[28611] + MEM[31195];
assign MEM[32598] = MEM[28612] + MEM[29379];
assign MEM[32599] = MEM[28613] + MEM[29010];
assign MEM[32600] = MEM[28614] + MEM[29892];
assign MEM[32601] = MEM[28615] + MEM[28841];
assign MEM[32602] = MEM[28618] + MEM[30254];
assign MEM[32603] = MEM[28622] + MEM[30442];
assign MEM[32604] = MEM[28627] + MEM[31718];
assign MEM[32605] = MEM[28628] + MEM[29858];
assign MEM[32606] = MEM[28630] + MEM[31250];
assign MEM[32607] = MEM[28631] + MEM[31294];
assign MEM[32608] = MEM[28633] + MEM[29796];
assign MEM[32609] = MEM[28634] + MEM[29767];
assign MEM[32610] = MEM[28640] + MEM[29323];
assign MEM[32611] = MEM[28641] + MEM[29319];
assign MEM[32612] = MEM[28644] + MEM[30438];
assign MEM[32613] = MEM[28646] + MEM[30774];
assign MEM[32614] = MEM[28648] + MEM[32068];
assign MEM[32615] = MEM[28649] + MEM[30759];
assign MEM[32616] = MEM[28652] + MEM[29365];
assign MEM[32617] = MEM[28653] + MEM[29327];
assign MEM[32618] = MEM[28655] + MEM[29469];
assign MEM[32619] = MEM[28656] + MEM[30681];
assign MEM[32620] = MEM[28657] + MEM[29539];
assign MEM[32621] = MEM[28664] + MEM[29933];
assign MEM[32622] = MEM[28666] + MEM[29357];
assign MEM[32623] = MEM[28667] + MEM[32039];
assign MEM[32624] = MEM[28668] + MEM[29550];
assign MEM[32625] = MEM[28669] + MEM[29364];
assign MEM[32626] = MEM[28673] + MEM[30009];
assign MEM[32627] = MEM[28674] + MEM[30092];
assign MEM[32628] = MEM[28680] + MEM[29998];
assign MEM[32629] = MEM[28681] + MEM[30076];
assign MEM[32630] = MEM[28682] + MEM[29074];
assign MEM[32631] = MEM[28684] + MEM[28881];
assign MEM[32632] = MEM[28687] + MEM[29149];
assign MEM[32633] = MEM[28688] + MEM[29462];
assign MEM[32634] = MEM[28691] + MEM[30709];
assign MEM[32635] = MEM[28693] + MEM[29741];
assign MEM[32636] = MEM[28694] + MEM[29812];
assign MEM[32637] = MEM[28695] + MEM[29649];
assign MEM[32638] = MEM[28697] + MEM[30536];
assign MEM[32639] = MEM[28698] + MEM[30995];
assign MEM[32640] = MEM[28699] + MEM[30197];
assign MEM[32641] = MEM[28700] + MEM[29446];
assign MEM[32642] = MEM[28702] + MEM[28807];
assign MEM[32643] = MEM[28703] + MEM[28836];
assign MEM[32644] = MEM[28705] + MEM[29143];
assign MEM[32645] = MEM[28713] + MEM[30175];
assign MEM[32646] = MEM[28714] + MEM[30630];
assign MEM[32647] = MEM[28716] + MEM[31064];
assign MEM[32648] = MEM[28723] + MEM[29300];
assign MEM[32649] = MEM[28726] + MEM[32050];
assign MEM[32650] = MEM[28729] + MEM[31451];
assign MEM[32651] = MEM[28731] + MEM[31649];
assign MEM[32652] = MEM[28732] + MEM[29460];
assign MEM[32653] = MEM[28736] + MEM[30309];
assign MEM[32654] = MEM[28737] + MEM[29508];
assign MEM[32655] = MEM[28741] + MEM[31612];
assign MEM[32656] = MEM[28745] + MEM[29823];
assign MEM[32657] = MEM[28746] + MEM[31855];
assign MEM[32658] = MEM[28748] + MEM[30094];
assign MEM[32659] = MEM[28749] + MEM[28932];
assign MEM[32660] = MEM[28750] + MEM[30136];
assign MEM[32661] = MEM[28751] + MEM[29564];
assign MEM[32662] = MEM[28755] + MEM[31989];
assign MEM[32663] = MEM[28756] + MEM[30859];
assign MEM[32664] = MEM[28759] + MEM[29224];
assign MEM[32665] = MEM[28760] + MEM[29809];
assign MEM[32666] = MEM[28761] + MEM[29162];
assign MEM[32667] = MEM[28765] + MEM[31296];
assign MEM[32668] = MEM[28767] + MEM[31114];
assign MEM[32669] = MEM[28768] + MEM[30727];
assign MEM[32670] = MEM[28769] + MEM[28904];
assign MEM[32671] = MEM[28770] + MEM[30218];
assign MEM[32672] = MEM[28772] + MEM[29474];
assign MEM[32673] = MEM[28775] + MEM[31080];
assign MEM[32674] = MEM[28777] + MEM[29737];
assign MEM[32675] = MEM[28779] + MEM[30029];
assign MEM[32676] = MEM[28785] + MEM[29900];
assign MEM[32677] = MEM[28786] + MEM[30070];
assign MEM[32678] = MEM[28788] + MEM[29360];
assign MEM[32679] = MEM[28789] + MEM[30731];
assign MEM[32680] = MEM[28791] + MEM[30604];
assign MEM[32681] = MEM[28796] + MEM[30974];
assign MEM[32682] = MEM[28801] + MEM[30538];
assign MEM[32683] = MEM[28802] + MEM[30396];
assign MEM[32684] = MEM[28805] + MEM[29131];
assign MEM[32685] = MEM[28808] + MEM[30758];
assign MEM[32686] = MEM[28811] + MEM[30374];
assign MEM[32687] = MEM[28812] + MEM[29778];
assign MEM[32688] = MEM[28816] + MEM[31892];
assign MEM[32689] = MEM[28821] + MEM[29620];
assign MEM[32690] = MEM[28822] + MEM[29363];
assign MEM[32691] = MEM[28824] + MEM[31719];
assign MEM[32692] = MEM[28828] + MEM[29618];
assign MEM[32693] = MEM[28830] + MEM[29376];
assign MEM[32694] = MEM[28832] + MEM[30751];
assign MEM[32695] = MEM[28833] + MEM[30702];
assign MEM[32696] = MEM[28835] + MEM[29921];
assign MEM[32697] = MEM[28837] + MEM[30496];
assign MEM[32698] = MEM[28838] + MEM[28864];
assign MEM[32699] = MEM[28839] + MEM[30384];
assign MEM[32700] = MEM[28840] + MEM[30967];
assign MEM[32701] = MEM[28842] + MEM[29494];
assign MEM[32702] = MEM[28846] + MEM[30434];
assign MEM[32703] = MEM[28849] + MEM[29167];
assign MEM[32704] = MEM[28850] + MEM[30036];
assign MEM[32705] = MEM[28852] + MEM[29994];
assign MEM[32706] = MEM[28854] + MEM[30337];
assign MEM[32707] = MEM[28856] + MEM[30924];
assign MEM[32708] = MEM[28857] + MEM[31100];
assign MEM[32709] = MEM[28860] + MEM[29247];
assign MEM[32710] = MEM[28861] + MEM[30730];
assign MEM[32711] = MEM[28867] + MEM[30541];
assign MEM[32712] = MEM[28869] + MEM[30863];
assign MEM[32713] = MEM[28871] + MEM[29366];
assign MEM[32714] = MEM[28873] + MEM[30500];
assign MEM[32715] = MEM[28875] + MEM[30649];
assign MEM[32716] = MEM[28876] + MEM[29960];
assign MEM[32717] = MEM[28877] + MEM[30880];
assign MEM[32718] = MEM[28878] + MEM[30260];
assign MEM[32719] = MEM[28879] + MEM[30628];
assign MEM[32720] = MEM[28880] + MEM[30295];
assign MEM[32721] = MEM[28882] + MEM[29316];
assign MEM[32722] = MEM[28884] + MEM[29075];
assign MEM[32723] = MEM[28887] + MEM[31007];
assign MEM[32724] = MEM[28889] + MEM[29752];
assign MEM[32725] = MEM[28891] + MEM[29771];
assign MEM[32726] = MEM[28894] + MEM[29486];
assign MEM[32727] = MEM[28897] + MEM[31227];
assign MEM[32728] = MEM[28898] + MEM[29166];
assign MEM[32729] = MEM[28900] + MEM[31117];
assign MEM[32730] = MEM[28905] + MEM[30525];
assign MEM[32731] = MEM[28907] + MEM[29711];
assign MEM[32732] = MEM[28909] + MEM[29108];
assign MEM[32733] = MEM[28911] + MEM[29047];
assign MEM[32734] = MEM[28914] + MEM[31392];
assign MEM[32735] = MEM[28915] + MEM[30741];
assign MEM[32736] = MEM[28916] + MEM[30571];
assign MEM[32737] = MEM[28917] + MEM[30552];
assign MEM[32738] = MEM[28920] + MEM[30146];
assign MEM[32739] = MEM[28921] + MEM[30835];
assign MEM[32740] = MEM[28922] + MEM[29296];
assign MEM[32741] = MEM[28925] + MEM[30674];
assign MEM[32742] = MEM[28928] + MEM[29385];
assign MEM[32743] = MEM[28931] + MEM[31428];
assign MEM[32744] = MEM[28937] + MEM[29160];
assign MEM[32745] = MEM[28938] + MEM[29217];
assign MEM[32746] = MEM[28939] + MEM[29259];
assign MEM[32747] = MEM[28941] + MEM[30382];
assign MEM[32748] = MEM[28942] + MEM[30444];
assign MEM[32749] = MEM[28943] + MEM[29787];
assign MEM[32750] = MEM[28945] + MEM[30133];
assign MEM[32751] = MEM[28947] + MEM[29342];
assign MEM[32752] = MEM[28949] + MEM[31665];
assign MEM[32753] = MEM[28950] + MEM[29712];
assign MEM[32754] = MEM[28951] + MEM[30237];
assign MEM[32755] = MEM[28954] + MEM[30847];
assign MEM[32756] = MEM[28955] + MEM[31405];
assign MEM[32757] = MEM[28957] + MEM[32106];
assign MEM[32758] = MEM[28961] + MEM[30342];
assign MEM[32759] = MEM[28962] + MEM[30851];
assign MEM[32760] = MEM[28966] + MEM[31016];
assign MEM[32761] = MEM[28968] + MEM[29936];
assign MEM[32762] = MEM[28970] + MEM[29838];
assign MEM[32763] = MEM[28971] + MEM[30929];
assign MEM[32764] = MEM[28976] + MEM[31008];
assign MEM[32765] = MEM[28977] + MEM[29887];
assign MEM[32766] = MEM[28978] + MEM[30306];
assign MEM[32767] = MEM[28980] + MEM[31097];
assign MEM[32768] = MEM[28981] + MEM[29860];
assign MEM[32769] = MEM[28986] + MEM[29635];
assign MEM[32770] = MEM[28988] + MEM[29703];
assign MEM[32771] = MEM[28992] + MEM[30728];
assign MEM[32772] = MEM[28993] + MEM[29488];
assign MEM[32773] = MEM[28994] + MEM[30334];
assign MEM[32774] = MEM[28996] + MEM[29170];
assign MEM[32775] = MEM[28997] + MEM[29558];
assign MEM[32776] = MEM[28998] + MEM[30931];
assign MEM[32777] = MEM[28999] + MEM[30307];
assign MEM[32778] = MEM[29000] + MEM[30243];
assign MEM[32779] = MEM[29002] + MEM[29263];
assign MEM[32780] = MEM[29003] + MEM[29230];
assign MEM[32781] = MEM[29004] + MEM[29671];
assign MEM[32782] = MEM[29005] + MEM[30498];
assign MEM[32783] = MEM[29006] + MEM[29980];
assign MEM[32784] = MEM[29008] + MEM[29485];
assign MEM[32785] = MEM[29009] + MEM[29358];
assign MEM[32786] = MEM[29014] + MEM[30348];
assign MEM[32787] = MEM[29015] + MEM[30310];
assign MEM[32788] = MEM[29016] + MEM[29690];
assign MEM[32789] = MEM[29017] + MEM[29732];
assign MEM[32790] = MEM[29018] + MEM[31236];
assign MEM[32791] = MEM[29020] + MEM[30058];
assign MEM[32792] = MEM[29024] + MEM[30166];
assign MEM[32793] = MEM[29025] + MEM[31124];
assign MEM[32794] = MEM[29026] + MEM[30869];
assign MEM[32795] = MEM[29027] + MEM[29456];
assign MEM[32796] = MEM[29030] + MEM[30071];
assign MEM[32797] = MEM[29034] + MEM[29148];
assign MEM[32798] = MEM[29037] + MEM[30471];
assign MEM[32799] = MEM[29038] + MEM[31166];
assign MEM[32800] = MEM[29039] + MEM[30723];
assign MEM[32801] = MEM[29041] + MEM[30028];
assign MEM[32802] = MEM[29044] + MEM[29299];
assign MEM[32803] = MEM[29049] + MEM[31073];
assign MEM[32804] = MEM[29051] + MEM[29696];
assign MEM[32805] = MEM[29052] + MEM[29877];
assign MEM[32806] = MEM[29054] + MEM[30117];
assign MEM[32807] = MEM[29055] + MEM[30823];
assign MEM[32808] = MEM[29056] + MEM[30431];
assign MEM[32809] = MEM[29057] + MEM[29262];
assign MEM[32810] = MEM[29064] + MEM[30497];
assign MEM[32811] = MEM[29066] + MEM[29653];
assign MEM[32812] = MEM[29068] + MEM[30796];
assign MEM[32813] = MEM[29070] + MEM[31631];
assign MEM[32814] = MEM[29071] + MEM[29808];
assign MEM[32815] = MEM[29073] + MEM[29229];
assign MEM[32816] = MEM[29076] + MEM[30683];
assign MEM[32817] = MEM[29077] + MEM[29626];
assign MEM[32818] = MEM[29078] + MEM[30079];
assign MEM[32819] = MEM[29081] + MEM[30779];
assign MEM[32820] = MEM[29082] + MEM[29610];
assign MEM[32821] = MEM[29083] + MEM[31365];
assign MEM[32822] = MEM[29085] + MEM[30679];
assign MEM[32823] = MEM[29087] + MEM[30208];
assign MEM[32824] = MEM[29089] + MEM[31182];
assign MEM[32825] = MEM[29090] + MEM[30477];
assign MEM[32826] = MEM[29091] + MEM[29305];
assign MEM[32827] = MEM[29092] + MEM[30128];
assign MEM[32828] = MEM[29093] + MEM[30129];
assign MEM[32829] = MEM[29094] + MEM[29422];
assign MEM[32830] = MEM[29095] + MEM[30816];
assign MEM[32831] = MEM[29096] + MEM[29806];
assign MEM[32832] = MEM[29098] + MEM[30145];
assign MEM[32833] = MEM[29099] + MEM[30399];
assign MEM[32834] = MEM[29100] + MEM[30032];
assign MEM[32835] = MEM[29102] + MEM[31464];
assign MEM[32836] = MEM[29103] + MEM[31871];
assign MEM[32837] = MEM[29104] + MEM[30909];
assign MEM[32838] = MEM[29106] + MEM[29890];
assign MEM[32839] = MEM[29107] + MEM[31988];
assign MEM[32840] = MEM[29109] + MEM[30961];
assign MEM[32841] = MEM[29111] + MEM[29280];
assign MEM[32842] = MEM[29113] + MEM[29307];
assign MEM[32843] = MEM[29115] + MEM[29594];
assign MEM[32844] = MEM[29117] + MEM[30209];
assign MEM[32845] = MEM[29120] + MEM[31506];
assign MEM[32846] = MEM[29122] + MEM[30242];
assign MEM[32847] = MEM[29127] + MEM[31038];
assign MEM[32848] = MEM[29128] + MEM[31148];
assign MEM[32849] = MEM[29132] + MEM[30614];
assign MEM[32850] = MEM[29136] + MEM[30357];
assign MEM[32851] = MEM[29138] + MEM[30775];
assign MEM[32852] = MEM[29139] + MEM[29962];
assign MEM[32853] = MEM[29140] + MEM[30879];
assign MEM[32854] = MEM[29145] + MEM[30824];
assign MEM[32855] = MEM[29147] + MEM[30921];
assign MEM[32856] = MEM[29150] + MEM[30400];
assign MEM[32857] = MEM[29154] + MEM[32322];
assign MEM[32858] = MEM[29159] + MEM[30177];
assign MEM[32859] = MEM[29161] + MEM[29941];
assign MEM[32860] = MEM[29163] + MEM[30566];
assign MEM[32861] = MEM[29165] + MEM[31002];
assign MEM[32862] = MEM[29169] + MEM[29467];
assign MEM[32863] = MEM[29173] + MEM[29315];
assign MEM[32864] = MEM[29177] + MEM[30225];
assign MEM[32865] = MEM[29181] + MEM[30417];
assign MEM[32866] = MEM[29185] + MEM[31961];
assign MEM[32867] = MEM[29188] + MEM[31116];
assign MEM[32868] = MEM[29193] + MEM[31449];
assign MEM[32869] = MEM[29197] + MEM[31229];
assign MEM[32870] = MEM[29200] + MEM[29995];
assign MEM[32871] = MEM[29201] + MEM[31386];
assign MEM[32872] = MEM[29203] + MEM[31371];
assign MEM[32873] = MEM[29205] + MEM[30113];
assign MEM[32874] = MEM[29207] + MEM[31135];
assign MEM[32875] = MEM[29209] + MEM[30724];
assign MEM[32876] = MEM[29210] + MEM[29672];
assign MEM[32877] = MEM[29212] + MEM[30427];
assign MEM[32878] = MEM[29213] + MEM[30600];
assign MEM[32879] = MEM[29218] + MEM[30221];
assign MEM[32880] = MEM[29220] + MEM[29851];
assign MEM[32881] = MEM[29221] + MEM[31489];
assign MEM[32882] = MEM[29223] + MEM[29384];
assign MEM[32883] = MEM[29225] + MEM[30805];
assign MEM[32884] = MEM[29226] + MEM[30047];
assign MEM[32885] = MEM[29227] + MEM[30726];
assign MEM[32886] = MEM[29232] + MEM[31280];
assign MEM[32887] = MEM[29233] + MEM[32396];
assign MEM[32888] = MEM[29235] + MEM[29616];
assign MEM[32889] = MEM[29237] + MEM[30229];
assign MEM[32890] = MEM[29240] + MEM[30335];
assign MEM[32891] = MEM[29242] + MEM[29546];
assign MEM[32892] = MEM[29245] + MEM[31085];
assign MEM[32893] = MEM[29246] + MEM[29527];
assign MEM[32894] = MEM[29248] + MEM[29837];
assign MEM[32895] = MEM[29250] + MEM[29830];
assign MEM[32896] = MEM[29253] + MEM[29770];
assign MEM[32897] = MEM[29254] + MEM[30349];
assign MEM[32898] = MEM[29255] + MEM[30772];
assign MEM[32899] = MEM[29256] + MEM[31933];
assign MEM[32900] = MEM[29258] + MEM[30663];
assign MEM[32901] = MEM[29260] + MEM[29502];
assign MEM[32902] = MEM[29261] + MEM[30543];
assign MEM[32903] = MEM[29266] + MEM[30697];
assign MEM[32904] = MEM[29272] + MEM[29479];
assign MEM[32905] = MEM[29273] + MEM[30200];
assign MEM[32906] = MEM[29274] + MEM[30352];
assign MEM[32907] = MEM[29276] + MEM[31686];
assign MEM[32908] = MEM[29277] + MEM[29832];
assign MEM[32909] = MEM[29278] + MEM[30275];
assign MEM[32910] = MEM[29283] + MEM[31717];
assign MEM[32911] = MEM[29284] + MEM[30096];
assign MEM[32912] = MEM[29287] + MEM[31336];
assign MEM[32913] = MEM[29288] + MEM[30168];
assign MEM[32914] = MEM[29291] + MEM[29563];
assign MEM[32915] = MEM[29293] + MEM[30783];
assign MEM[32916] = MEM[29294] + MEM[30919];
assign MEM[32917] = MEM[29295] + MEM[31150];
assign MEM[32918] = MEM[29297] + MEM[30052];
assign MEM[32919] = MEM[29301] + MEM[30794];
assign MEM[32920] = MEM[29306] + MEM[29440];
assign MEM[32921] = MEM[29309] + MEM[29430];
assign MEM[32922] = MEM[29313] + MEM[31233];
assign MEM[32923] = MEM[29314] + MEM[29940];
assign MEM[32924] = MEM[29317] + MEM[30188];
assign MEM[32925] = MEM[29318] + MEM[29785];
assign MEM[32926] = MEM[29320] + MEM[30170];
assign MEM[32927] = MEM[29321] + MEM[30401];
assign MEM[32928] = MEM[29322] + MEM[31217];
assign MEM[32929] = MEM[29328] + MEM[30239];
assign MEM[32930] = MEM[29330] + MEM[30110];
assign MEM[32931] = MEM[29332] + MEM[30888];
assign MEM[32932] = MEM[29335] + MEM[31487];
assign MEM[32933] = MEM[29336] + MEM[31448];
assign MEM[32934] = MEM[29337] + MEM[30786];
assign MEM[32935] = MEM[29338] + MEM[30652];
assign MEM[32936] = MEM[29339] + MEM[29810];
assign MEM[32937] = MEM[29341] + MEM[31325];
assign MEM[32938] = MEM[29345] + MEM[30285];
assign MEM[32939] = MEM[29351] + MEM[30872];
assign MEM[32940] = MEM[29352] + MEM[31643];
assign MEM[32941] = MEM[29353] + MEM[30472];
assign MEM[32942] = MEM[29355] + MEM[30296];
assign MEM[32943] = MEM[29356] + MEM[29782];
assign MEM[32944] = MEM[29361] + MEM[29856];
assign MEM[32945] = MEM[29367] + MEM[31032];
assign MEM[32946] = MEM[29369] + MEM[31264];
assign MEM[32947] = MEM[29371] + MEM[29878];
assign MEM[32948] = MEM[29373] + MEM[29917];
assign MEM[32949] = MEM[29374] + MEM[29648];
assign MEM[32950] = MEM[29377] + MEM[30761];
assign MEM[32951] = MEM[29378] + MEM[30998];
assign MEM[32952] = MEM[29382] + MEM[30433];
assign MEM[32953] = MEM[29383] + MEM[29819];
assign MEM[32954] = MEM[29387] + MEM[30426];
assign MEM[32955] = MEM[29388] + MEM[31446];
assign MEM[32956] = MEM[29389] + MEM[30176];
assign MEM[32957] = MEM[29390] + MEM[32264];
assign MEM[32958] = MEM[29394] + MEM[29604];
assign MEM[32959] = MEM[29395] + MEM[30699];
assign MEM[32960] = MEM[29396] + MEM[32330];
assign MEM[32961] = MEM[29397] + MEM[29595];
assign MEM[32962] = MEM[29398] + MEM[30403];
assign MEM[32963] = MEM[29399] + MEM[29911];
assign MEM[32964] = MEM[29401] + MEM[31318];
assign MEM[32965] = MEM[29403] + MEM[30535];
assign MEM[32966] = MEM[29404] + MEM[29896];
assign MEM[32967] = MEM[29405] + MEM[32103];
assign MEM[32968] = MEM[29406] + MEM[30347];
assign MEM[32969] = MEM[29409] + MEM[31543];
assign MEM[32970] = MEM[29411] + MEM[31591];
assign MEM[32971] = MEM[29415] + MEM[29772];
assign MEM[32972] = MEM[29417] + MEM[30682];
assign MEM[32973] = MEM[29421] + MEM[31492];
assign MEM[32974] = MEM[29423] + MEM[31323];
assign MEM[32975] = MEM[29424] + MEM[31054];
assign MEM[32976] = MEM[29426] + MEM[30523];
assign MEM[32977] = MEM[29428] + MEM[30388];
assign MEM[32978] = MEM[29429] + MEM[32037];
assign MEM[32979] = MEM[29433] + MEM[30184];
assign MEM[32980] = MEM[29434] + MEM[31082];
assign MEM[32981] = MEM[29436] + MEM[30707];
assign MEM[32982] = MEM[29437] + MEM[30018];
assign MEM[32983] = MEM[29438] + MEM[29891];
assign MEM[32984] = MEM[29441] + MEM[30559];
assign MEM[32985] = MEM[29442] + MEM[31526];
assign MEM[32986] = MEM[29444] + MEM[32055];
assign MEM[32987] = MEM[29445] + MEM[30279];
assign MEM[32988] = MEM[29447] + MEM[30091];
assign MEM[32989] = MEM[29449] + MEM[29768];
assign MEM[32990] = MEM[29450] + MEM[30986];
assign MEM[32991] = MEM[29451] + MEM[29817];
assign MEM[32992] = MEM[29452] + MEM[30095];
assign MEM[32993] = MEM[29455] + MEM[31340];
assign MEM[32994] = MEM[29463] + MEM[30005];
assign MEM[32995] = MEM[29465] + MEM[29499];
assign MEM[32996] = MEM[29471] + MEM[30840];
assign MEM[32997] = MEM[29473] + MEM[31027];
assign MEM[32998] = MEM[29475] + MEM[30488];
assign MEM[32999] = MEM[29476] + MEM[31216];
assign MEM[33000] = MEM[29478] + MEM[31121];
assign MEM[33001] = MEM[29482] + MEM[30395];
assign MEM[33002] = MEM[29483] + MEM[29742];
assign MEM[33003] = MEM[29489] + MEM[30629];
assign MEM[33004] = MEM[29490] + MEM[29735];
assign MEM[33005] = MEM[29491] + MEM[30084];
assign MEM[33006] = MEM[29493] + MEM[31720];
assign MEM[33007] = MEM[29495] + MEM[30641];
assign MEM[33008] = MEM[29498] + MEM[31103];
assign MEM[33009] = MEM[29500] + MEM[30875];
assign MEM[33010] = MEM[29503] + MEM[30769];
assign MEM[33011] = MEM[29504] + MEM[30620];
assign MEM[33012] = MEM[29507] + MEM[31573];
assign MEM[33013] = MEM[29510] + MEM[30361];
assign MEM[33014] = MEM[29513] + MEM[31426];
assign MEM[33015] = MEM[29518] + MEM[29598];
assign MEM[33016] = MEM[29532] + MEM[30623];
assign MEM[33017] = MEM[29533] + MEM[31888];
assign MEM[33018] = MEM[29534] + MEM[29942];
assign MEM[33019] = MEM[29535] + MEM[31138];
assign MEM[33020] = MEM[29536] + MEM[30885];
assign MEM[33021] = MEM[29545] + MEM[29766];
assign MEM[33022] = MEM[29547] + MEM[30321];
assign MEM[33023] = MEM[29548] + MEM[32409];
assign MEM[33024] = MEM[29549] + MEM[31224];
assign MEM[33025] = MEM[29551] + MEM[29996];
assign MEM[33026] = MEM[29552] + MEM[29920];
assign MEM[33027] = MEM[29556] + MEM[31026];
assign MEM[33028] = MEM[29559] + MEM[32478];
assign MEM[33029] = MEM[29561] + MEM[30428];
assign MEM[33030] = MEM[29562] + MEM[32245];
assign MEM[33031] = MEM[29566] + MEM[31397];
assign MEM[33032] = MEM[29567] + MEM[30464];
assign MEM[33033] = MEM[29568] + MEM[30481];
assign MEM[33034] = MEM[29569] + MEM[29855];
assign MEM[33035] = MEM[29570] + MEM[29882];
assign MEM[33036] = MEM[29571] + MEM[31049];
assign MEM[33037] = MEM[29573] + MEM[29985];
assign MEM[33038] = MEM[29575] + MEM[30276];
assign MEM[33039] = MEM[29576] + MEM[30367];
assign MEM[33040] = MEM[29580] + MEM[31067];
assign MEM[33041] = MEM[29582] + MEM[30037];
assign MEM[33042] = MEM[29583] + MEM[30745];
assign MEM[33043] = MEM[29584] + MEM[30778];
assign MEM[33044] = MEM[29586] + MEM[30913];
assign MEM[33045] = MEM[29590] + MEM[29749];
assign MEM[33046] = MEM[29591] + MEM[30414];
assign MEM[33047] = MEM[29593] + MEM[30643];
assign MEM[33048] = MEM[29597] + MEM[31088];
assign MEM[33049] = MEM[29599] + MEM[31158];
assign MEM[33050] = MEM[29600] + MEM[31516];
assign MEM[33051] = MEM[29602] + MEM[30920];
assign MEM[33052] = MEM[29603] + MEM[31347];
assign MEM[33053] = MEM[29608] + MEM[30033];
assign MEM[33054] = MEM[29612] + MEM[31646];
assign MEM[33055] = MEM[29613] + MEM[30518];
assign MEM[33056] = MEM[29614] + MEM[30404];
assign MEM[33057] = MEM[29615] + MEM[31929];
assign MEM[33058] = MEM[29622] + MEM[31495];
assign MEM[33059] = MEM[29624] + MEM[31128];
assign MEM[33060] = MEM[29625] + MEM[30125];
assign MEM[33061] = MEM[29628] + MEM[31161];
assign MEM[33062] = MEM[29630] + MEM[29814];
assign MEM[33063] = MEM[29631] + MEM[29979];
assign MEM[33064] = MEM[29633] + MEM[30547];
assign MEM[33065] = MEM[29636] + MEM[30292];
assign MEM[33066] = MEM[29638] + MEM[31075];
assign MEM[33067] = MEM[29641] + MEM[31101];
assign MEM[33068] = MEM[29644] + MEM[30645];
assign MEM[33069] = MEM[29646] + MEM[31880];
assign MEM[33070] = MEM[29650] + MEM[30150];
assign MEM[33071] = MEM[29651] + MEM[30943];
assign MEM[33072] = MEM[29656] + MEM[31439];
assign MEM[33073] = MEM[29657] + MEM[32152];
assign MEM[33074] = MEM[29659] + MEM[30561];
assign MEM[33075] = MEM[29660] + MEM[30003];
assign MEM[33076] = MEM[29662] + MEM[30189];
assign MEM[33077] = MEM[29664] + MEM[31163];
assign MEM[33078] = MEM[29666] + MEM[31382];
assign MEM[33079] = MEM[29667] + MEM[30676];
assign MEM[33080] = MEM[29669] + MEM[32334];
assign MEM[33081] = MEM[29670] + MEM[31728];
assign MEM[33082] = MEM[29673] + MEM[31076];
assign MEM[33083] = MEM[29674] + MEM[30385];
assign MEM[33084] = MEM[29675] + MEM[30550];
assign MEM[33085] = MEM[29676] + MEM[31307];
assign MEM[33086] = MEM[29678] + MEM[30680];
assign MEM[33087] = MEM[29680] + MEM[30114];
assign MEM[33088] = MEM[29681] + MEM[30733];
assign MEM[33089] = MEM[29682] + MEM[31193];
assign MEM[33090] = MEM[29684] + MEM[30540];
assign MEM[33091] = MEM[29686] + MEM[30486];
assign MEM[33092] = MEM[29687] + MEM[31132];
assign MEM[33093] = MEM[29689] + MEM[30960];
assign MEM[33094] = MEM[29691] + MEM[30735];
assign MEM[33095] = MEM[29692] + MEM[31122];
assign MEM[33096] = MEM[29693] + MEM[31313];
assign MEM[33097] = MEM[29695] + MEM[31154];
assign MEM[33098] = MEM[29697] + MEM[31019];
assign MEM[33099] = MEM[29700] + MEM[31208];
assign MEM[33100] = MEM[29702] + MEM[31519];
assign MEM[33101] = MEM[29705] + MEM[31772];
assign MEM[33102] = MEM[29706] + MEM[30320];
assign MEM[33103] = MEM[29709] + MEM[32118];
assign MEM[33104] = MEM[29716] + MEM[32376];
assign MEM[33105] = MEM[29717] + MEM[32826];
assign MEM[33106] = MEM[29718] + MEM[31493];
assign MEM[33107] = MEM[29724] + MEM[32648];
assign MEM[33108] = MEM[29725] + MEM[31180];
assign MEM[33109] = MEM[29728] + MEM[32167];
assign MEM[33110] = MEM[29731] + MEM[31206];
assign MEM[33111] = MEM[29738] + MEM[32412];
assign MEM[33112] = MEM[29739] + MEM[31355];
assign MEM[33113] = MEM[29740] + MEM[32510];
assign MEM[33114] = MEM[29743] + MEM[31510];
assign MEM[33115] = MEM[29744] + MEM[31266];
assign MEM[33116] = MEM[29746] + MEM[31984];
assign MEM[33117] = MEM[29751] + MEM[30817];
assign MEM[33118] = MEM[29755] + MEM[30976];
assign MEM[33119] = MEM[29756] + MEM[32125];
assign MEM[33120] = MEM[29759] + MEM[31339];
assign MEM[33121] = MEM[29760] + MEM[30088];
assign MEM[33122] = MEM[29769] + MEM[31857];
assign MEM[33123] = MEM[29775] + MEM[31587];
assign MEM[33124] = MEM[29776] + MEM[32161];
assign MEM[33125] = MEM[29779] + MEM[31574];
assign MEM[33126] = MEM[29781] + MEM[32098];
assign MEM[33127] = MEM[29783] + MEM[32159];
assign MEM[33128] = MEM[29795] + MEM[32262];
assign MEM[33129] = MEM[29799] + MEM[32020];
assign MEM[33130] = MEM[29800] + MEM[32598];
assign MEM[33131] = MEM[29803] + MEM[32099];
assign MEM[33132] = MEM[29804] + MEM[30989];
assign MEM[33133] = MEM[29805] + MEM[32056];
assign MEM[33134] = MEM[29807] + MEM[31260];
assign MEM[33135] = MEM[29813] + MEM[31477];
assign MEM[33136] = MEM[29815] + MEM[31239];
assign MEM[33137] = MEM[29818] + MEM[31832];
assign MEM[33138] = MEM[29820] + MEM[31671];
assign MEM[33139] = MEM[29822] + MEM[31955];
assign MEM[33140] = MEM[29824] + MEM[32258];
assign MEM[33141] = MEM[29826] + MEM[31674];
assign MEM[33142] = MEM[29827] + MEM[31104];
assign MEM[33143] = MEM[29828] + MEM[31035];
assign MEM[33144] = MEM[29831] + MEM[31647];
assign MEM[33145] = MEM[29833] + MEM[32538];
assign MEM[33146] = MEM[29834] + MEM[32429];
assign MEM[33147] = MEM[29836] + MEM[30789];
assign MEM[33148] = MEM[29840] + MEM[31262];
assign MEM[33149] = MEM[29842] + MEM[31808];
assign MEM[33150] = MEM[29844] + MEM[31560];
assign MEM[33151] = MEM[29845] + MEM[32449];
assign MEM[33152] = MEM[29846] + MEM[31848];
assign MEM[33153] = MEM[29848] + MEM[31839];
assign MEM[33154] = MEM[29853] + MEM[31762];
assign MEM[33155] = MEM[29854] + MEM[30752];
assign MEM[33156] = MEM[29861] + MEM[31376];
assign MEM[33157] = MEM[29862] + MEM[31462];
assign MEM[33158] = MEM[29863] + MEM[31828];
assign MEM[33159] = MEM[29871] + MEM[31583];
assign MEM[33160] = MEM[29872] + MEM[31727];
assign MEM[33161] = MEM[29875] + MEM[31454];
assign MEM[33162] = MEM[29879] + MEM[31308];
assign MEM[33163] = MEM[29880] + MEM[31185];
assign MEM[33164] = MEM[29883] + MEM[30753];
assign MEM[33165] = MEM[29893] + MEM[31678];
assign MEM[33166] = MEM[29894] + MEM[31242];
assign MEM[33167] = MEM[29897] + MEM[32348];
assign MEM[33168] = MEM[29898] + MEM[31069];
assign MEM[33169] = MEM[29899] + MEM[31090];
assign MEM[33170] = MEM[29901] + MEM[31442];
assign MEM[33171] = MEM[29904] + MEM[32362];
assign MEM[33172] = MEM[29906] + MEM[31902];
assign MEM[33173] = MEM[29907] + MEM[32361];
assign MEM[33174] = MEM[29908] + MEM[32678];
assign MEM[33175] = MEM[29910] + MEM[31901];
assign MEM[33176] = MEM[29912] + MEM[32289];
assign MEM[33177] = MEM[29915] + MEM[30368];
assign MEM[33178] = MEM[29916] + MEM[32841];
assign MEM[33179] = MEM[29918] + MEM[32301];
assign MEM[33180] = MEM[29919] + MEM[31981];
assign MEM[33181] = MEM[29922] + MEM[31079];
assign MEM[33182] = MEM[29926] + MEM[31249];
assign MEM[33183] = MEM[29944] + MEM[32172];
assign MEM[33184] = MEM[29949] + MEM[32433];
assign MEM[33185] = MEM[29953] + MEM[31589];
assign MEM[33186] = MEM[29957] + MEM[31691];
assign MEM[33187] = MEM[29958] + MEM[32137];
assign MEM[33188] = MEM[29961] + MEM[31126];
assign MEM[33189] = MEM[29964] + MEM[31432];
assign MEM[33190] = MEM[29970] + MEM[32326];
assign MEM[33191] = MEM[29975] + MEM[31326];
assign MEM[33192] = MEM[29976] + MEM[31406];
assign MEM[33193] = MEM[29977] + MEM[32207];
assign MEM[33194] = MEM[29981] + MEM[31542];
assign MEM[33195] = MEM[29983] + MEM[31134];
assign MEM[33196] = MEM[29986] + MEM[32625];
assign MEM[33197] = MEM[29988] + MEM[31884];
assign MEM[33198] = MEM[29989] + MEM[31547];
assign MEM[33199] = MEM[29992] + MEM[32036];
assign MEM[33200] = MEM[29997] + MEM[31197];
assign MEM[33201] = MEM[30001] + MEM[31570];
assign MEM[33202] = MEM[30010] + MEM[31805];
assign MEM[33203] = MEM[30012] + MEM[31044];
assign MEM[33204] = MEM[30014] + MEM[32033];
assign MEM[33205] = MEM[30015] + MEM[30390];
assign MEM[33206] = MEM[30016] + MEM[31697];
assign MEM[33207] = MEM[30017] + MEM[32426];
assign MEM[33208] = MEM[30023] + MEM[31967];
assign MEM[33209] = MEM[30024] + MEM[30814];
assign MEM[33210] = MEM[30026] + MEM[31730];
assign MEM[33211] = MEM[30030] + MEM[31734];
assign MEM[33212] = MEM[30031] + MEM[31771];
assign MEM[33213] = MEM[30035] + MEM[31541];
assign MEM[33214] = MEM[30038] + MEM[32028];
assign MEM[33215] = MEM[30039] + MEM[31115];
assign MEM[33216] = MEM[30040] + MEM[31960];
assign MEM[33217] = MEM[30042] + MEM[31342];
assign MEM[33218] = MEM[30044] + MEM[31780];
assign MEM[33219] = MEM[30048] + MEM[31928];
assign MEM[33220] = MEM[30051] + MEM[31680];
assign MEM[33221] = MEM[30054] + MEM[32503];
assign MEM[33222] = MEM[30055] + MEM[31982];
assign MEM[33223] = MEM[30056] + MEM[31877];
assign MEM[33224] = MEM[30059] + MEM[30954];
assign MEM[33225] = MEM[30062] + MEM[31363];
assign MEM[33226] = MEM[30063] + MEM[31757];
assign MEM[33227] = MEM[30064] + MEM[30811];
assign MEM[33228] = MEM[30066] + MEM[31247];
assign MEM[33229] = MEM[30067] + MEM[32809];
assign MEM[33230] = MEM[30068] + MEM[30820];
assign MEM[33231] = MEM[30077] + MEM[31463];
assign MEM[33232] = MEM[30081] + MEM[31230];
assign MEM[33233] = MEM[30083] + MEM[32456];
assign MEM[33234] = MEM[30086] + MEM[32862];
assign MEM[33235] = MEM[30087] + MEM[31020];
assign MEM[33236] = MEM[30089] + MEM[32795];
assign MEM[33237] = MEM[30090] + MEM[31952];
assign MEM[33238] = MEM[30098] + MEM[32029];
assign MEM[33239] = MEM[30102] + MEM[31231];
assign MEM[33240] = MEM[30103] + MEM[32690];
assign MEM[33241] = MEM[30104] + MEM[31765];
assign MEM[33242] = MEM[30105] + MEM[32785];
assign MEM[33243] = MEM[30107] + MEM[31200];
assign MEM[33244] = MEM[30111] + MEM[31838];
assign MEM[33245] = MEM[30118] + MEM[31240];
assign MEM[33246] = MEM[30123] + MEM[31751];
assign MEM[33247] = MEM[30124] + MEM[31913];
assign MEM[33248] = MEM[30127] + MEM[31438];
assign MEM[33249] = MEM[30130] + MEM[31858];
assign MEM[33250] = MEM[30131] + MEM[31530];
assign MEM[33251] = MEM[30134] + MEM[31941];
assign MEM[33252] = MEM[30135] + MEM[31990];
assign MEM[33253] = MEM[30140] + MEM[32312];
assign MEM[33254] = MEM[30142] + MEM[33005];
assign MEM[33255] = MEM[30147] + MEM[31859];
assign MEM[33256] = MEM[30149] + MEM[31275];
assign MEM[33257] = MEM[30153] + MEM[31424];
assign MEM[33258] = MEM[30155] + MEM[32529];
assign MEM[33259] = MEM[30157] + MEM[31750];
assign MEM[33260] = MEM[30163] + MEM[32643];
assign MEM[33261] = MEM[30167] + MEM[31679];
assign MEM[33262] = MEM[30173] + MEM[32008];
assign MEM[33263] = MEM[30174] + MEM[31501];
assign MEM[33264] = MEM[30178] + MEM[32077];
assign MEM[33265] = MEM[30179] + MEM[31940];
assign MEM[33266] = MEM[30182] + MEM[32246];
assign MEM[33267] = MEM[30185] + MEM[31498];
assign MEM[33268] = MEM[30191] + MEM[31466];
assign MEM[33269] = MEM[30193] + MEM[31557];
assign MEM[33270] = MEM[30194] + MEM[32057];
assign MEM[33271] = MEM[30195] + MEM[31975];
assign MEM[33272] = MEM[30196] + MEM[31087];
assign MEM[33273] = MEM[30201] + MEM[32904];
assign MEM[33274] = MEM[30202] + MEM[31974];
assign MEM[33275] = MEM[30211] + MEM[32296];
assign MEM[33276] = MEM[30212] + MEM[31947];
assign MEM[33277] = MEM[30213] + MEM[31287];
assign MEM[33278] = MEM[30216] + MEM[31891];
assign MEM[33279] = MEM[30222] + MEM[31258];
assign MEM[33280] = MEM[30224] + MEM[31830];
assign MEM[33281] = MEM[30228] + MEM[31301];
assign MEM[33282] = MEM[30230] + MEM[30837];
assign MEM[33283] = MEM[30232] + MEM[31253];
assign MEM[33284] = MEM[30233] + MEM[31630];
assign MEM[33285] = MEM[30241] + MEM[31849];
assign MEM[33286] = MEM[30244] + MEM[31531];
assign MEM[33287] = MEM[30248] + MEM[32366];
assign MEM[33288] = MEM[30252] + MEM[31559];
assign MEM[33289] = MEM[30255] + MEM[31171];
assign MEM[33290] = MEM[30257] + MEM[32155];
assign MEM[33291] = MEM[30261] + MEM[31496];
assign MEM[33292] = MEM[30264] + MEM[32590];
assign MEM[33293] = MEM[30268] + MEM[32481];
assign MEM[33294] = MEM[30272] + MEM[32219];
assign MEM[33295] = MEM[30274] + MEM[31306];
assign MEM[33296] = MEM[30282] + MEM[32428];
assign MEM[33297] = MEM[30283] + MEM[31851];
assign MEM[33298] = MEM[30289] + MEM[32368];
assign MEM[33299] = MEM[30293] + MEM[31726];
assign MEM[33300] = MEM[30297] + MEM[31351];
assign MEM[33301] = MEM[30300] + MEM[31458];
assign MEM[33302] = MEM[30302] + MEM[30827];
assign MEM[33303] = MEM[30303] + MEM[31759];
assign MEM[33304] = MEM[30305] + MEM[31912];
assign MEM[33305] = MEM[30316] + MEM[31806];
assign MEM[33306] = MEM[30323] + MEM[31070];
assign MEM[33307] = MEM[30324] + MEM[31532];
assign MEM[33308] = MEM[30326] + MEM[32303];
assign MEM[33309] = MEM[30327] + MEM[32274];
assign MEM[33310] = MEM[30336] + MEM[32591];
assign MEM[33311] = MEM[30340] + MEM[31962];
assign MEM[33312] = MEM[30344] + MEM[31648];
assign MEM[33313] = MEM[30354] + MEM[32522];
assign MEM[33314] = MEM[30355] + MEM[32599];
assign MEM[33315] = MEM[30358] + MEM[31181];
assign MEM[33316] = MEM[30363] + MEM[31914];
assign MEM[33317] = MEM[30364] + MEM[32102];
assign MEM[33318] = MEM[30366] + MEM[32035];
assign MEM[33319] = MEM[30373] + MEM[31846];
assign MEM[33320] = MEM[30375] + MEM[31710];
assign MEM[33321] = MEM[30379] + MEM[32592];
assign MEM[33322] = MEM[30386] + MEM[32047];
assign MEM[33323] = MEM[30391] + MEM[31165];
assign MEM[33324] = MEM[30397] + MEM[31349];
assign MEM[33325] = MEM[30407] + MEM[32000];
assign MEM[33326] = MEM[30408] + MEM[32147];
assign MEM[33327] = MEM[30410] + MEM[32052];
assign MEM[33328] = MEM[30415] + MEM[31919];
assign MEM[33329] = MEM[30418] + MEM[32224];
assign MEM[33330] = MEM[30421] + MEM[32624];
assign MEM[33331] = MEM[30424] + MEM[32270];
assign MEM[33332] = MEM[30429] + MEM[31825];
assign MEM[33333] = MEM[30430] + MEM[32129];
assign MEM[33334] = MEM[30437] + MEM[32797];
assign MEM[33335] = MEM[30443] + MEM[31983];
assign MEM[33336] = MEM[30445] + MEM[31517];
assign MEM[33337] = MEM[30451] + MEM[31580];
assign MEM[33338] = MEM[30453] + MEM[32005];
assign MEM[33339] = MEM[30454] + MEM[32064];
assign MEM[33340] = MEM[30455] + MEM[32622];
assign MEM[33341] = MEM[30456] + MEM[32183];
assign MEM[33342] = MEM[30458] + MEM[31729];
assign MEM[33343] = MEM[30461] + MEM[31797];
assign MEM[33344] = MEM[30466] + MEM[32530];
assign MEM[33345] = MEM[30469] + MEM[31317];
assign MEM[33346] = MEM[30474] + MEM[31659];
assign MEM[33347] = MEM[30476] + MEM[32065];
assign MEM[33348] = MEM[30478] + MEM[31595];
assign MEM[33349] = MEM[30479] + MEM[31092];
assign MEM[33350] = MEM[30487] + MEM[32024];
assign MEM[33351] = MEM[30491] + MEM[31977];
assign MEM[33352] = MEM[30492] + MEM[31434];
assign MEM[33353] = MEM[30495] + MEM[31670];
assign MEM[33354] = MEM[30501] + MEM[32081];
assign MEM[33355] = MEM[30502] + MEM[31611];
assign MEM[33356] = MEM[30503] + MEM[32504];
assign MEM[33357] = MEM[30507] + MEM[31698];
assign MEM[33358] = MEM[30508] + MEM[31567];
assign MEM[33359] = MEM[30509] + MEM[32382];
assign MEM[33360] = MEM[30511] + MEM[31309];
assign MEM[33361] = MEM[30514] + MEM[31869];
assign MEM[33362] = MEM[30517] + MEM[32038];
assign MEM[33363] = MEM[30519] + MEM[31895];
assign MEM[33364] = MEM[30520] + MEM[32022];
assign MEM[33365] = MEM[30521] + MEM[31137];
assign MEM[33366] = MEM[30522] + MEM[31485];
assign MEM[33367] = MEM[30524] + MEM[32373];
assign MEM[33368] = MEM[30530] + MEM[31110];
assign MEM[33369] = MEM[30539] + MEM[31943];
assign MEM[33370] = MEM[30542] + MEM[31508];
assign MEM[33371] = MEM[30544] + MEM[32482];
assign MEM[33372] = MEM[30546] + MEM[31337];
assign MEM[33373] = MEM[30557] + MEM[32358];
assign MEM[33374] = MEM[30560] + MEM[31390];
assign MEM[33375] = MEM[30562] + MEM[32631];
assign MEM[33376] = MEM[30563] + MEM[31436];
assign MEM[33377] = MEM[30564] + MEM[31875];
assign MEM[33378] = MEM[30570] + MEM[31421];
assign MEM[33379] = MEM[30573] + MEM[32091];
assign MEM[33380] = MEM[30576] + MEM[32189];
assign MEM[33381] = MEM[30579] + MEM[32239];
assign MEM[33382] = MEM[30581] + MEM[32512];
assign MEM[33383] = MEM[30587] + MEM[32143];
assign MEM[33384] = MEM[30589] + MEM[32435];
assign MEM[33385] = MEM[30590] + MEM[32944];
assign MEM[33386] = MEM[30591] + MEM[31948];
assign MEM[33387] = MEM[30592] + MEM[32413];
assign MEM[33388] = MEM[30594] + MEM[32009];
assign MEM[33389] = MEM[30597] + MEM[32498];
assign MEM[33390] = MEM[30598] + MEM[32774];
assign MEM[33391] = MEM[30599] + MEM[32444];
assign MEM[33392] = MEM[30603] + MEM[32046];
assign MEM[33393] = MEM[30607] + MEM[31297];
assign MEM[33394] = MEM[30608] + MEM[31764];
assign MEM[33395] = MEM[30609] + MEM[31059];
assign MEM[33396] = MEM[30615] + MEM[31699];
assign MEM[33397] = MEM[30616] + MEM[31608];
assign MEM[33398] = MEM[30619] + MEM[32532];
assign MEM[33399] = MEM[30621] + MEM[32582];
assign MEM[33400] = MEM[30626] + MEM[32323];
assign MEM[33401] = MEM[30632] + MEM[32437];
assign MEM[33402] = MEM[30636] + MEM[32784];
assign MEM[33403] = MEM[30638] + MEM[31894];
assign MEM[33404] = MEM[30639] + MEM[31430];
assign MEM[33405] = MEM[30644] + MEM[31978];
assign MEM[33406] = MEM[30646] + MEM[31700];
assign MEM[33407] = MEM[30647] + MEM[31636];
assign MEM[33408] = MEM[30651] + MEM[31125];
assign MEM[33409] = MEM[30653] + MEM[31702];
assign MEM[33410] = MEM[30654] + MEM[31835];
assign MEM[33411] = MEM[30655] + MEM[31601];
assign MEM[33412] = MEM[30656] + MEM[32130];
assign MEM[33413] = MEM[30659] + MEM[32013];
assign MEM[33414] = MEM[30660] + MEM[31744];
assign MEM[33415] = MEM[30662] + MEM[31521];
assign MEM[33416] = MEM[30669] + MEM[32703];
assign MEM[33417] = MEM[30673] + MEM[32215];
assign MEM[33418] = MEM[30678] + MEM[32048];
assign MEM[33419] = MEM[30685] + MEM[31470];
assign MEM[33420] = MEM[30689] + MEM[31709];
assign MEM[33421] = MEM[30690] + MEM[31372];
assign MEM[33422] = MEM[30694] + MEM[31707];
assign MEM[33423] = MEM[30703] + MEM[31527];
assign MEM[33424] = MEM[30705] + MEM[32117];
assign MEM[33425] = MEM[30706] + MEM[31904];
assign MEM[33426] = MEM[30711] + MEM[31528];
assign MEM[33427] = MEM[30713] + MEM[32108];
assign MEM[33428] = MEM[30714] + MEM[31922];
assign MEM[33429] = MEM[30717] + MEM[32181];
assign MEM[33430] = MEM[30719] + MEM[32051];
assign MEM[33431] = MEM[30721] + MEM[31136];
assign MEM[33432] = MEM[30722] + MEM[32772];
assign MEM[33433] = MEM[30738] + MEM[32399];
assign MEM[33434] = MEM[30739] + MEM[31118];
assign MEM[33435] = MEM[30742] + MEM[32133];
assign MEM[33436] = MEM[30744] + MEM[31809];
assign MEM[33437] = MEM[30748] + MEM[31754];
assign MEM[33438] = MEM[30750] + MEM[32463];
assign MEM[33439] = MEM[30757] + MEM[31415];
assign MEM[33440] = MEM[30764] + MEM[32165];
assign MEM[33441] = MEM[30766] + MEM[31656];
assign MEM[33442] = MEM[30767] + MEM[32356];
assign MEM[33443] = MEM[30771] + MEM[31949];
assign MEM[33444] = MEM[30777] + MEM[31844];
assign MEM[33445] = MEM[30780] + MEM[32006];
assign MEM[33446] = MEM[30782] + MEM[31548];
assign MEM[33447] = MEM[30785] + MEM[31860];
assign MEM[33448] = MEM[30792] + MEM[32288];
assign MEM[33449] = MEM[30793] + MEM[31733];
assign MEM[33450] = MEM[30798] + MEM[32438];
assign MEM[33451] = MEM[30799] + MEM[32726];
assign MEM[33452] = MEM[30802] + MEM[32032];
assign MEM[33453] = MEM[30806] + MEM[31388];
assign MEM[33454] = MEM[30807] + MEM[32462];
assign MEM[33455] = MEM[30808] + MEM[31921];
assign MEM[33456] = MEM[30815] + MEM[31916];
assign MEM[33457] = MEM[30822] + MEM[31711];
assign MEM[33458] = MEM[30828] + MEM[31964];
assign MEM[33459] = MEM[30831] + MEM[31576];
assign MEM[33460] = MEM[30832] + MEM[31621];
assign MEM[33461] = MEM[30836] + MEM[32484];
assign MEM[33462] = MEM[30842] + MEM[32260];
assign MEM[33463] = MEM[30848] + MEM[31712];
assign MEM[33464] = MEM[30853] + MEM[31481];
assign MEM[33465] = MEM[30854] + MEM[31514];
assign MEM[33466] = MEM[30855] + MEM[32017];
assign MEM[33467] = MEM[30858] + MEM[32421];
assign MEM[33468] = MEM[30860] + MEM[32265];
assign MEM[33469] = MEM[30861] + MEM[32417];
assign MEM[33470] = MEM[30862] + MEM[31915];
assign MEM[33471] = MEM[30865] + MEM[31781];
assign MEM[33472] = MEM[30871] + MEM[32223];
assign MEM[33473] = MEM[30873] + MEM[31786];
assign MEM[33474] = MEM[30876] + MEM[31564];
assign MEM[33475] = MEM[30886] + MEM[32333];
assign MEM[33476] = MEM[30890] + MEM[31556];
assign MEM[33477] = MEM[30892] + MEM[31803];
assign MEM[33478] = MEM[30893] + MEM[32448];
assign MEM[33479] = MEM[30897] + MEM[31684];
assign MEM[33480] = MEM[30898] + MEM[31578];
assign MEM[33481] = MEM[30899] + MEM[31333];
assign MEM[33482] = MEM[30901] + MEM[32187];
assign MEM[33483] = MEM[30903] + MEM[31893];
assign MEM[33484] = MEM[30904] + MEM[31954];
assign MEM[33485] = MEM[30906] + MEM[32151];
assign MEM[33486] = MEM[30910] + MEM[32287];
assign MEM[33487] = MEM[30911] + MEM[32594];
assign MEM[33488] = MEM[30912] + MEM[32175];
assign MEM[33489] = MEM[30914] + MEM[32318];
assign MEM[33490] = MEM[30916] + MEM[31605];
assign MEM[33491] = MEM[30918] + MEM[32814];
assign MEM[33492] = MEM[30922] + MEM[31735];
assign MEM[33493] = MEM[30925] + MEM[32618];
assign MEM[33494] = MEM[30934] + MEM[32882];
assign MEM[33495] = MEM[30936] + MEM[31742];
assign MEM[33496] = MEM[30944] + MEM[31474];
assign MEM[33497] = MEM[30946] + MEM[32015];
assign MEM[33498] = MEM[30948] + MEM[31833];
assign MEM[33499] = MEM[30950] + MEM[32163];
assign MEM[33500] = MEM[30953] + MEM[32231];
assign MEM[33501] = MEM[30956] + MEM[31865];
assign MEM[33502] = MEM[30963] + MEM[32491];
assign MEM[33503] = MEM[30964] + MEM[32441];
assign MEM[33504] = MEM[30965] + MEM[32460];
assign MEM[33505] = MEM[30970] + MEM[32222];
assign MEM[33506] = MEM[30972] + MEM[32012];
assign MEM[33507] = MEM[30973] + MEM[31932];
assign MEM[33508] = MEM[30975] + MEM[32141];
assign MEM[33509] = MEM[30980] + MEM[32476];
assign MEM[33510] = MEM[30982] + MEM[31886];
assign MEM[33511] = MEM[30984] + MEM[32418];
assign MEM[33512] = MEM[30988] + MEM[32178];
assign MEM[33513] = MEM[30992] + MEM[31628];
assign MEM[33514] = MEM[30993] + MEM[32042];
assign MEM[33515] = MEM[30994] + MEM[32578];
assign MEM[33516] = MEM[30996] + MEM[32025];
assign MEM[33517] = MEM[31000] + MEM[32104];
assign MEM[33518] = MEM[31004] + MEM[32011];
assign MEM[33519] = MEM[31005] + MEM[32401];
assign MEM[33520] = MEM[31010] + MEM[32938];
assign MEM[33521] = MEM[31012] + MEM[32629];
assign MEM[33522] = MEM[31013] + MEM[32218];
assign MEM[33523] = MEM[31015] + MEM[32567];
assign MEM[33524] = MEM[31021] + MEM[32393];
assign MEM[33525] = MEM[31025] + MEM[32229];
assign MEM[33526] = MEM[31031] + MEM[32390];
assign MEM[33527] = MEM[31034] + MEM[31739];
assign MEM[33528] = MEM[31036] + MEM[32226];
assign MEM[33529] = MEM[31037] + MEM[32263];
assign MEM[33530] = MEM[31040] + MEM[32779];
assign MEM[33531] = MEM[31041] + MEM[32466];
assign MEM[33532] = MEM[31043] + MEM[31873];
assign MEM[33533] = MEM[31047] + MEM[32442];
assign MEM[33534] = MEM[31051] + MEM[31937];
assign MEM[33535] = MEM[31052] + MEM[32721];
assign MEM[33536] = MEM[31053] + MEM[32953];
assign MEM[33537] = MEM[31055] + MEM[32929];
assign MEM[33538] = MEM[31058] + MEM[32641];
assign MEM[33539] = MEM[31062] + MEM[32234];
assign MEM[33540] = MEM[31065] + MEM[32588];
assign MEM[33541] = MEM[31068] + MEM[32403];
assign MEM[33542] = MEM[31072] + MEM[32256];
assign MEM[33543] = MEM[31077] + MEM[32605];
assign MEM[33544] = MEM[31081] + MEM[32352];
assign MEM[33545] = MEM[31086] + MEM[32235];
assign MEM[33546] = MEM[31091] + MEM[32436];
assign MEM[33547] = MEM[31093] + MEM[31968];
assign MEM[33548] = MEM[31096] + MEM[32633];
assign MEM[33549] = MEM[31099] + MEM[33021];
assign MEM[33550] = MEM[31102] + MEM[31768];
assign MEM[33551] = MEM[31105] + MEM[32526];
assign MEM[33552] = MEM[31109] + MEM[32420];
assign MEM[33553] = MEM[31123] + MEM[31845];
assign MEM[33554] = MEM[31130] + MEM[31994];
assign MEM[33555] = MEM[31133] + MEM[32683];
assign MEM[33556] = MEM[31140] + MEM[32134];
assign MEM[33557] = MEM[31142] + MEM[32063];
assign MEM[33558] = MEM[31143] + MEM[32562];
assign MEM[33559] = MEM[31152] + MEM[31898];
assign MEM[33560] = MEM[31155] + MEM[32394];
assign MEM[33561] = MEM[31156] + MEM[32286];
assign MEM[33562] = MEM[31162] + MEM[32744];
assign MEM[33563] = MEM[31167] + MEM[32030];
assign MEM[33564] = MEM[31168] + MEM[32897];
assign MEM[33565] = MEM[31169] + MEM[33015];
assign MEM[33566] = MEM[31172] + MEM[32549];
assign MEM[33567] = MEM[31178] + MEM[32573];
assign MEM[33568] = MEM[31179] + MEM[32071];
assign MEM[33569] = MEM[31190] + MEM[32781];
assign MEM[33570] = MEM[31191] + MEM[31931];
assign MEM[33571] = MEM[31192] + MEM[32295];
assign MEM[33572] = MEM[31194] + MEM[32320];
assign MEM[33573] = MEM[31198] + MEM[31936];
assign MEM[33574] = MEM[31201] + MEM[31522];
assign MEM[33575] = MEM[31202] + MEM[32812];
assign MEM[33576] = MEM[31204] + MEM[32736];
assign MEM[33577] = MEM[31211] + MEM[32116];
assign MEM[33578] = MEM[31215] + MEM[32961];
assign MEM[33579] = MEM[31218] + MEM[32440];
assign MEM[33580] = MEM[31219] + MEM[32268];
assign MEM[33581] = MEM[31222] + MEM[32305];
assign MEM[33582] = MEM[31232] + MEM[31625];
assign MEM[33583] = MEM[31241] + MEM[31864];
assign MEM[33584] = MEM[31243] + MEM[32948];
assign MEM[33585] = MEM[31255] + MEM[32539];
assign MEM[33586] = MEM[31256] + MEM[32253];
assign MEM[33587] = MEM[31257] + MEM[32656];
assign MEM[33588] = MEM[31268] + MEM[32921];
assign MEM[33589] = MEM[31272] + MEM[32010];
assign MEM[33590] = MEM[31273] + MEM[32676];
assign MEM[33591] = MEM[31274] + MEM[32045];
assign MEM[33592] = MEM[31282] + MEM[32855];
assign MEM[33593] = MEM[31286] + MEM[32346];
assign MEM[33594] = MEM[31292] + MEM[32820];
assign MEM[33595] = MEM[31295] + MEM[32644];
assign MEM[33596] = MEM[31298] + MEM[32121];
assign MEM[33597] = MEM[31300] + MEM[32873];
assign MEM[33598] = MEM[31302] + MEM[32095];
assign MEM[33599] = MEM[31310] + MEM[32389];
assign MEM[33600] = MEM[31312] + MEM[32076];
assign MEM[33601] = MEM[31314] + MEM[31867];
assign MEM[33602] = MEM[31315] + MEM[32715];
assign MEM[33603] = MEM[31316] + MEM[32559];
assign MEM[33604] = MEM[31319] + MEM[32331];
assign MEM[33605] = MEM[31320] + MEM[32551];
assign MEM[33606] = MEM[31321] + MEM[33025];
assign MEM[33607] = MEM[31322] + MEM[32865];
assign MEM[33608] = MEM[31328] + MEM[32319];
assign MEM[33609] = MEM[31330] + MEM[32019];
assign MEM[33610] = MEM[31332] + MEM[32164];
assign MEM[33611] = MEM[31338] + MEM[33102];
assign MEM[33612] = MEM[31346] + MEM[32082];
assign MEM[33613] = MEM[31352] + MEM[32459];
assign MEM[33614] = MEM[31358] + MEM[32293];
assign MEM[33615] = MEM[31361] + MEM[32817];
assign MEM[33616] = MEM[31366] + MEM[32423];
assign MEM[33617] = MEM[31368] + MEM[32828];
assign MEM[33618] = MEM[31370] + MEM[32609];
assign MEM[33619] = MEM[31377] + MEM[32672];
assign MEM[33620] = MEM[31380] + MEM[31675];
assign MEM[33621] = MEM[31381] + MEM[32146];
assign MEM[33622] = MEM[31387] + MEM[32771];
assign MEM[33623] = MEM[31395] + MEM[32843];
assign MEM[33624] = MEM[31396] + MEM[32901];
assign MEM[33625] = MEM[31398] + MEM[33094];
assign MEM[33626] = MEM[31399] + MEM[31824];
assign MEM[33627] = MEM[31401] + MEM[32994];
assign MEM[33628] = MEM[31402] + MEM[32351];
assign MEM[33629] = MEM[31408] + MEM[32859];
assign MEM[33630] = MEM[31410] + MEM[32365];
assign MEM[33631] = MEM[31414] + MEM[32205];
assign MEM[33632] = MEM[31422] + MEM[32699];
assign MEM[33633] = MEM[31427] + MEM[32652];
assign MEM[33634] = MEM[31433] + MEM[31694];
assign MEM[33635] = MEM[31443] + MEM[32898];
assign MEM[33636] = MEM[31445] + MEM[32976];
assign MEM[33637] = MEM[31450] + MEM[32513];
assign MEM[33638] = MEM[31455] + MEM[32596];
assign MEM[33639] = MEM[31461] + MEM[32314];
assign MEM[33640] = MEM[31465] + MEM[32492];
assign MEM[33641] = MEM[31467] + MEM[31966];
assign MEM[33642] = MEM[31472] + MEM[32124];
assign MEM[33643] = MEM[31473] + MEM[32391];
assign MEM[33644] = MEM[31476] + MEM[32770];
assign MEM[33645] = MEM[31480] + MEM[31993];
assign MEM[33646] = MEM[31482] + MEM[32555];
assign MEM[33647] = MEM[31486] + MEM[32272];
assign MEM[33648] = MEM[31488] + MEM[32294];
assign MEM[33649] = MEM[31491] + MEM[32834];
assign MEM[33650] = MEM[31502] + MEM[32706];
assign MEM[33651] = MEM[31503] + MEM[32925];
assign MEM[33652] = MEM[31505] + MEM[32619];
assign MEM[33653] = MEM[31507] + MEM[32328];
assign MEM[33654] = MEM[31509] + MEM[32354];
assign MEM[33655] = MEM[31512] + MEM[32233];
assign MEM[33656] = MEM[31513] + MEM[32515];
assign MEM[33657] = MEM[31515] + MEM[32664];
assign MEM[33658] = MEM[31518] + MEM[33095];
assign MEM[33659] = MEM[31523] + MEM[32544];
assign MEM[33660] = MEM[31533] + MEM[32431];
assign MEM[33661] = MEM[31535] + MEM[32364];
assign MEM[33662] = MEM[31540] + MEM[32796];
assign MEM[33663] = MEM[31553] + MEM[32769];
assign MEM[33664] = MEM[31555] + MEM[33065];
assign MEM[33665] = MEM[31558] + MEM[32693];
assign MEM[33666] = MEM[31561] + MEM[32156];
assign MEM[33667] = MEM[31566] + MEM[32569];
assign MEM[33668] = MEM[31569] + MEM[32406];
assign MEM[33669] = MEM[31571] + MEM[32684];
assign MEM[33670] = MEM[31575] + MEM[32507];
assign MEM[33671] = MEM[31577] + MEM[32838];
assign MEM[33672] = MEM[31579] + MEM[32891];
assign MEM[33673] = MEM[31582] + MEM[32202];
assign MEM[33674] = MEM[31585] + MEM[32004];
assign MEM[33675] = MEM[31592] + MEM[33046];
assign MEM[33676] = MEM[31598] + MEM[32278];
assign MEM[33677] = MEM[31603] + MEM[32031];
assign MEM[33678] = MEM[31604] + MEM[32827];
assign MEM[33679] = MEM[31606] + MEM[32864];
assign MEM[33680] = MEM[31615] + MEM[32833];
assign MEM[33681] = MEM[31618] + MEM[31792];
assign MEM[33682] = MEM[31622] + MEM[32930];
assign MEM[33683] = MEM[31623] + MEM[32892];
assign MEM[33684] = MEM[31624] + MEM[32475];
assign MEM[33685] = MEM[31626] + MEM[32811];
assign MEM[33686] = MEM[31629] + MEM[32560];
assign MEM[33687] = MEM[31632] + MEM[32877];
assign MEM[33688] = MEM[31635] + MEM[32991];
assign MEM[33689] = MEM[31639] + MEM[33002];
assign MEM[33690] = MEM[31640] + MEM[32724];
assign MEM[33691] = MEM[31652] + MEM[32908];
assign MEM[33692] = MEM[31653] + MEM[32277];
assign MEM[33693] = MEM[31654] + MEM[32638];
assign MEM[33694] = MEM[31658] + MEM[32720];
assign MEM[33695] = MEM[31661] + MEM[32489];
assign MEM[33696] = MEM[31677] + MEM[32616];
assign MEM[33697] = MEM[31682] + MEM[32924];
assign MEM[33698] = MEM[31687] + MEM[32696];
assign MEM[33699] = MEM[31688] + MEM[32170];
assign MEM[33700] = MEM[31689] + MEM[32537];
assign MEM[33701] = MEM[31690] + MEM[32708];
assign MEM[33702] = MEM[31693] + MEM[32452];
assign MEM[33703] = MEM[31695] + MEM[32627];
assign MEM[33704] = MEM[31696] + MEM[32485];
assign MEM[33705] = MEM[31705] + MEM[32284];
assign MEM[33706] = MEM[31708] + MEM[33142];
assign MEM[33707] = MEM[31737] + MEM[32850];
assign MEM[33708] = MEM[31741] + MEM[33032];
assign MEM[33709] = MEM[31743] + MEM[32842];
assign MEM[33710] = MEM[31745] + MEM[32608];
assign MEM[33711] = MEM[31748] + MEM[32837];
assign MEM[33712] = MEM[31755] + MEM[32640];
assign MEM[33713] = MEM[31763] + MEM[32816];
assign MEM[33714] = MEM[31766] + MEM[32249];
assign MEM[33715] = MEM[31767] + MEM[32992];
assign MEM[33716] = MEM[31769] + MEM[32153];
assign MEM[33717] = MEM[31773] + MEM[32832];
assign MEM[33718] = MEM[31776] + MEM[32761];
assign MEM[33719] = MEM[31779] + MEM[32470];
assign MEM[33720] = MEM[31790] + MEM[32439];
assign MEM[33721] = MEM[31795] + MEM[32210];
assign MEM[33722] = MEM[31799] + MEM[32801];
assign MEM[33723] = MEM[31800] + MEM[32411];
assign MEM[33724] = MEM[31804] + MEM[32177];
assign MEM[33725] = MEM[31813] + MEM[32791];
assign MEM[33726] = MEM[31817] + MEM[32603];
assign MEM[33727] = MEM[31818] + MEM[32981];
assign MEM[33728] = MEM[31821] + MEM[32917];
assign MEM[33729] = MEM[31836] + MEM[32963];
assign MEM[33730] = MEM[31840] + MEM[32502];
assign MEM[33731] = MEM[31842] + MEM[32765];
assign MEM[33732] = MEM[31847] + MEM[32653];
assign MEM[33733] = MEM[31850] + MEM[32600];
assign MEM[33734] = MEM[31853] + MEM[32639];
assign MEM[33735] = MEM[31854] + MEM[32909];
assign MEM[33736] = MEM[31856] + MEM[32751];
assign MEM[33737] = MEM[31868] + MEM[32692];
assign MEM[33738] = MEM[31870] + MEM[33074];
assign MEM[33739] = MEM[31872] + MEM[32360];
assign MEM[33740] = MEM[31874] + MEM[32941];
assign MEM[33741] = MEM[31878] + MEM[32645];
assign MEM[33742] = MEM[31879] + MEM[32499];
assign MEM[33743] = MEM[31899] + MEM[33121];
assign MEM[33744] = MEM[31903] + MEM[32325];
assign MEM[33745] = MEM[31907] + MEM[32902];
assign MEM[33746] = MEM[31908] + MEM[32990];
assign MEM[33747] = MEM[31911] + MEM[32982];
assign MEM[33748] = MEM[31917] + MEM[33134];
assign MEM[33749] = MEM[31918] + MEM[32807];
assign MEM[33750] = MEM[31923] + MEM[32918];
assign MEM[33751] = MEM[31924] + MEM[32145];
assign MEM[33752] = MEM[31925] + MEM[32988];
assign MEM[33753] = MEM[31926] + MEM[33041];
assign MEM[33754] = MEM[31938] + MEM[32942];
assign MEM[33755] = MEM[31945] + MEM[32329];
assign MEM[33756] = MEM[31946] + MEM[32875];
assign MEM[33757] = MEM[31953] + MEM[33415];
assign MEM[33758] = MEM[31956] + MEM[32900];
assign MEM[33759] = MEM[31963] + MEM[32822];
assign MEM[33760] = MEM[31969] + MEM[33163];
assign MEM[33761] = MEM[31973] + MEM[32896];
assign MEM[33762] = MEM[31979] + MEM[32800];
assign MEM[33763] = MEM[31987] + MEM[32472];
assign MEM[33764] = MEM[31992] + MEM[32890];
assign MEM[33765] = MEM[31996] + MEM[32705];
assign MEM[33766] = MEM[32002] + MEM[32716];
assign MEM[33767] = MEM[32023] + MEM[32977];
assign MEM[33768] = MEM[32026] + MEM[33365];
assign MEM[33769] = MEM[32053] + MEM[33035];
assign MEM[33770] = MEM[32060] + MEM[32554];
assign MEM[33771] = MEM[32061] + MEM[33421];
assign MEM[33772] = MEM[32069] + MEM[33099];
assign MEM[33773] = MEM[32074] + MEM[32686];
assign MEM[33774] = MEM[32083] + MEM[32553];
assign MEM[33775] = MEM[32084] + MEM[33089];
assign MEM[33776] = MEM[32086] + MEM[32753];
assign MEM[33777] = MEM[32093] + MEM[33083];
assign MEM[33778] = MEM[32094] + MEM[32749];
assign MEM[33779] = MEM[32097] + MEM[32636];
assign MEM[33780] = MEM[32100] + MEM[32840];
assign MEM[33781] = MEM[32110] + MEM[32670];
assign MEM[33782] = MEM[32111] + MEM[32762];
assign MEM[33783] = MEM[32112] + MEM[33257];
assign MEM[33784] = MEM[32113] + MEM[32725];
assign MEM[33785] = MEM[32119] + MEM[33052];
assign MEM[33786] = MEM[32120] + MEM[32488];
assign MEM[33787] = MEM[32122] + MEM[32867];
assign MEM[33788] = MEM[32126] + MEM[33090];
assign MEM[33789] = MEM[32127] + MEM[32665];
assign MEM[33790] = MEM[32128] + MEM[32806];
assign MEM[33791] = MEM[32144] + MEM[32985];
assign MEM[33792] = MEM[32148] + MEM[33239];
assign MEM[33793] = MEM[32150] + MEM[32913];
assign MEM[33794] = MEM[32160] + MEM[32970];
assign MEM[33795] = MEM[32162] + MEM[33047];
assign MEM[33796] = MEM[32168] + MEM[32928];
assign MEM[33797] = MEM[32169] + MEM[32767];
assign MEM[33798] = MEM[32173] + MEM[32956];
assign MEM[33799] = MEM[32174] + MEM[33210];
assign MEM[33800] = MEM[32179] + MEM[33185];
assign MEM[33801] = MEM[32184] + MEM[33031];
assign MEM[33802] = MEM[32193] + MEM[32773];
assign MEM[33803] = MEM[32194] + MEM[33426];
assign MEM[33804] = MEM[32195] + MEM[32974];
assign MEM[33805] = MEM[32199] + MEM[33209];
assign MEM[33806] = MEM[32201] + MEM[33282];
assign MEM[33807] = MEM[32203] + MEM[32758];
assign MEM[33808] = MEM[32206] + MEM[33053];
assign MEM[33809] = MEM[32209] + MEM[32695];
assign MEM[33810] = MEM[32211] + MEM[32714];
assign MEM[33811] = MEM[32213] + MEM[33376];
assign MEM[33812] = MEM[32216] + MEM[32818];
assign MEM[33813] = MEM[32217] + MEM[33056];
assign MEM[33814] = MEM[32225] + MEM[33059];
assign MEM[33815] = MEM[32227] + MEM[33169];
assign MEM[33816] = MEM[32228] + MEM[32525];
assign MEM[33817] = MEM[32230] + MEM[32747];
assign MEM[33818] = MEM[32240] + MEM[33345];
assign MEM[33819] = MEM[32255] + MEM[32989];
assign MEM[33820] = MEM[32257] + MEM[32858];
assign MEM[33821] = MEM[32267] + MEM[33369];
assign MEM[33822] = MEM[32275] + MEM[33004];
assign MEM[33823] = MEM[32276] + MEM[33681];
assign MEM[33824] = MEM[32279] + MEM[33199];
assign MEM[33825] = MEM[32280] + MEM[32783];
assign MEM[33826] = MEM[32281] + MEM[32979];
assign MEM[33827] = MEM[32290] + MEM[32969];
assign MEM[33828] = MEM[32291] + MEM[33040];
assign MEM[33829] = MEM[32292] + MEM[33091];
assign MEM[33830] = MEM[32299] + MEM[33123];
assign MEM[33831] = MEM[32300] + MEM[32455];
assign MEM[33832] = MEM[32316] + MEM[32876];
assign MEM[33833] = MEM[32332] + MEM[32935];
assign MEM[33834] = MEM[32339] + MEM[32884];
assign MEM[33835] = MEM[32341] + MEM[33003];
assign MEM[33836] = MEM[32342] + MEM[33036];
assign MEM[33837] = MEM[32349] + MEM[32894];
assign MEM[33838] = MEM[32374] + MEM[32968];
assign MEM[33839] = MEM[32377] + MEM[33001];
assign MEM[33840] = MEM[32378] + MEM[32748];
assign MEM[33841] = MEM[32380] + MEM[32848];
assign MEM[33842] = MEM[32384] + MEM[32906];
assign MEM[33843] = MEM[32387] + MEM[33414];
assign MEM[33844] = MEM[32407] + MEM[33100];
assign MEM[33845] = MEM[32414] + MEM[33039];
assign MEM[33846] = MEM[32430] + MEM[33204];
assign MEM[33847] = MEM[32447] + MEM[33349];
assign MEM[33848] = MEM[32451] + MEM[33038];
assign MEM[33849] = MEM[32457] + MEM[33447];
assign MEM[33850] = MEM[32468] + MEM[33228];
assign MEM[33851] = MEM[32471] + MEM[33474];
assign MEM[33852] = MEM[32477] + MEM[32793];
assign MEM[33853] = MEM[32509] + MEM[33194];
assign MEM[33854] = MEM[32518] + MEM[33591];
assign MEM[33855] = MEM[32520] + MEM[32746];
assign MEM[33856] = MEM[32541] + MEM[32794];
assign MEM[33857] = MEM[32543] + MEM[33136];
assign MEM[33858] = MEM[32546] + MEM[33168];
assign MEM[33859] = MEM[32550] + MEM[33499];
assign MEM[33860] = MEM[32563] + MEM[33235];
assign MEM[33861] = MEM[32568] + MEM[33195];
assign MEM[33862] = MEM[32574] + MEM[33319];
assign MEM[33863] = MEM[32581] + MEM[33550];
assign MEM[33864] = MEM[32584] + MEM[33599];
assign MEM[33865] = MEM[32587] + MEM[32803];
assign MEM[33866] = MEM[32595] + MEM[32825];
assign MEM[33867] = MEM[32601] + MEM[33197];
assign MEM[33868] = MEM[32610] + MEM[33404];
assign MEM[33869] = MEM[32611] + MEM[33328];
assign MEM[33870] = MEM[32617] + MEM[33252];
assign MEM[33871] = MEM[32620] + MEM[33180];
assign MEM[33872] = MEM[32630] + MEM[33397];
assign MEM[33873] = MEM[32632] + MEM[33686];
assign MEM[33874] = MEM[32634] + MEM[33598];
assign MEM[33875] = MEM[32637] + MEM[33427];
assign MEM[33876] = MEM[32642] + MEM[33076];
assign MEM[33877] = MEM[32659] + MEM[33058];
assign MEM[33878] = MEM[32661] + MEM[33085];
assign MEM[33879] = MEM[32689] + MEM[33531];
assign MEM[33880] = MEM[32698] + MEM[33490];
assign MEM[33881] = MEM[32701] + MEM[33113];
assign MEM[33882] = MEM[32704] + MEM[33645];
assign MEM[33883] = MEM[32709] + MEM[33306];
assign MEM[33884] = MEM[32722] + MEM[32910];
assign MEM[33885] = MEM[32728] + MEM[33051];
assign MEM[33886] = MEM[32732] + MEM[33612];
assign MEM[33887] = MEM[32740] + MEM[33342];
assign MEM[33888] = MEM[32742] + MEM[33372];
assign MEM[33889] = MEM[32745] + MEM[33000];
assign MEM[33890] = MEM[32775] + MEM[33283];
assign MEM[33891] = MEM[32780] + MEM[33389];
assign MEM[33892] = MEM[32788] + MEM[33222];
assign MEM[33893] = MEM[32792] + MEM[33462];
assign MEM[33894] = MEM[32802] + MEM[33106];
assign MEM[33895] = MEM[32804] + MEM[33563];
assign MEM[33896] = MEM[32815] + MEM[33013];
assign MEM[33897] = MEM[32829] + MEM[33301];
assign MEM[33898] = MEM[32863] + MEM[33454];
assign MEM[33899] = MEM[32880] + MEM[33512];
assign MEM[33900] = MEM[32888] + MEM[33470];
assign MEM[33901] = MEM[32893] + MEM[33303];
assign MEM[33902] = MEM[32914] + MEM[33151];
assign MEM[33903] = MEM[32920] + MEM[33542];
assign MEM[33904] = MEM[32949] + MEM[33483];
assign MEM[33905] = MEM[32958] + MEM[33524];
assign MEM[33906] = MEM[32971] + MEM[33553];
assign MEM[33907] = MEM[32995] + MEM[33191];
assign MEM[33908] = MEM[33029] + MEM[33533];
assign MEM[33909] = MEM[33033] + MEM[33626];
assign MEM[33910] = MEM[33034] + MEM[33660];
assign MEM[33911] = MEM[33045] + MEM[33657];
assign MEM[33912] = MEM[33060] + MEM[33476];
assign MEM[33913] = MEM[33071] + MEM[33855];
assign MEM[33914] = MEM[33075] + MEM[33573];
assign MEM[33915] = MEM[33098] + MEM[33730];
assign MEM[33916] = MEM[33155] + MEM[33736];
assign MEM[33917] = MEM[33227] + MEM[33574];
assign MEM[33918] = MEM[33243] + MEM[33696];
assign MEM[33919] = MEM[5] + MEM[542];
assign MEM[33920] = MEM[7] + MEM[70];
assign MEM[33921] = MEM[13] + MEM[46];
assign MEM[33922] = MEM[15] + MEM[303];
assign MEM[33923] = MEM[21] + MEM[95];
assign MEM[33924] = MEM[22] + MEM[380];
assign MEM[33925] = MEM[38] + MEM[270];
assign MEM[33926] = MEM[45] + MEM[78];
assign MEM[33927] = MEM[54] + MEM[415];
assign MEM[33928] = MEM[61] + MEM[255];
assign MEM[33929] = MEM[71] + MEM[359];
assign MEM[33930] = MEM[79] + MEM[183];
assign MEM[33931] = MEM[93] + MEM[411];
assign MEM[33932] = MEM[94] + MEM[901];
assign MEM[33933] = MEM[110] + MEM[262];
assign MEM[33934] = MEM[117] + MEM[175];
assign MEM[33935] = MEM[119] + MEM[661];
assign MEM[33936] = MEM[133] + MEM[570];
assign MEM[33937] = MEM[134] + MEM[269];
assign MEM[33938] = MEM[135] + MEM[213];
assign MEM[33939] = MEM[143] + MEM[751];
assign MEM[33940] = MEM[158] + MEM[529];
assign MEM[33941] = MEM[165] + MEM[354];
assign MEM[33942] = MEM[167] + MEM[316];
assign MEM[33943] = MEM[181] + MEM[239];
assign MEM[33944] = MEM[182] + MEM[522];
assign MEM[33945] = MEM[190] + MEM[293];
assign MEM[33946] = MEM[205] + MEM[557];
assign MEM[33947] = MEM[221] + MEM[930];
assign MEM[33948] = MEM[222] + MEM[310];
assign MEM[33949] = MEM[223] + MEM[455];
assign MEM[33950] = MEM[237] + MEM[758];
assign MEM[33951] = MEM[238] + MEM[759];
assign MEM[33952] = MEM[277] + MEM[862];
assign MEM[33953] = MEM[284] + MEM[746];
assign MEM[33954] = MEM[292] + MEM[747];
assign MEM[33955] = MEM[294] + MEM[322];
assign MEM[33956] = MEM[295] + MEM[338];
assign MEM[33957] = MEM[306] + MEM[530];
assign MEM[33958] = MEM[315] + MEM[373];
assign MEM[33959] = MEM[318] + MEM[603];
assign MEM[33960] = MEM[319] + MEM[386];
assign MEM[33961] = MEM[323] + MEM[540];
assign MEM[33962] = MEM[339] + MEM[850];
assign MEM[33963] = MEM[347] + MEM[1091];
assign MEM[33964] = MEM[350] + MEM[583];
assign MEM[33965] = MEM[358] + MEM[679];
assign MEM[33966] = MEM[363] + MEM[514];
assign MEM[33967] = MEM[365] + MEM[585];
assign MEM[33968] = MEM[367] + MEM[547];
assign MEM[33969] = MEM[370] + MEM[395];
assign MEM[33970] = MEM[371] + MEM[382];
assign MEM[33971] = MEM[378] + MEM[389];
assign MEM[33972] = MEM[379] + MEM[952];
assign MEM[33973] = MEM[381] + MEM[728];
assign MEM[33974] = MEM[383] + MEM[517];
assign MEM[33975] = MEM[399] + MEM[516];
assign MEM[33976] = MEM[422] + MEM[493];
assign MEM[33977] = MEM[423] + MEM[781];
assign MEM[33978] = MEM[438] + MEM[470];
assign MEM[33979] = MEM[471] + MEM[709];
assign MEM[33980] = MEM[483] + MEM[727];
assign MEM[33981] = MEM[487] + MEM[771];
assign MEM[33982] = MEM[503] + MEM[662];
assign MEM[33983] = MEM[510] + MEM[551];
assign MEM[33984] = MEM[511] + MEM[655];
assign MEM[33985] = MEM[518] + MEM[846];
assign MEM[33986] = MEM[534] + MEM[733];
assign MEM[33987] = MEM[545] + MEM[579];
assign MEM[33988] = MEM[558] + MEM[604];
assign MEM[33989] = MEM[559] + MEM[834];
assign MEM[33990] = MEM[561] + MEM[692];
assign MEM[33991] = MEM[562] + MEM[566];
assign MEM[33992] = MEM[564] + MEM[590];
assign MEM[33993] = MEM[573] + MEM[992];
assign MEM[33994] = MEM[586] + MEM[601];
assign MEM[33995] = MEM[593] + MEM[1487];
assign MEM[33996] = MEM[598] + MEM[1442];
assign MEM[33997] = MEM[599] + MEM[610];
assign MEM[33998] = MEM[602] + MEM[677];
assign MEM[33999] = MEM[607] + MEM[693];
assign MEM[34000] = MEM[619] + MEM[1079];
assign MEM[34001] = MEM[627] + MEM[927];
assign MEM[34002] = MEM[628] + MEM[756];
assign MEM[34003] = MEM[635] + MEM[685];
assign MEM[34004] = MEM[644] + MEM[950];
assign MEM[34005] = MEM[646] + MEM[722];
assign MEM[34006] = MEM[652] + MEM[822];
assign MEM[34007] = MEM[663] + MEM[813];
assign MEM[34008] = MEM[686] + MEM[1141];
assign MEM[34009] = MEM[695] + MEM[940];
assign MEM[34010] = MEM[711] + MEM[744];
assign MEM[34011] = MEM[719] + MEM[740];
assign MEM[34012] = MEM[730] + MEM[937];
assign MEM[34013] = MEM[741] + MEM[876];
assign MEM[34014] = MEM[748] + MEM[773];
assign MEM[34015] = MEM[749] + MEM[999];
assign MEM[34016] = MEM[757] + MEM[811];
assign MEM[34017] = MEM[760] + MEM[789];
assign MEM[34018] = MEM[766] + MEM[1510];
assign MEM[34019] = MEM[769] + MEM[919];
assign MEM[34020] = MEM[772] + MEM[1030];
assign MEM[34021] = MEM[779] + MEM[838];
assign MEM[34022] = MEM[790] + MEM[797];
assign MEM[34023] = MEM[794] + MEM[852];
assign MEM[34024] = MEM[805] + MEM[1076];
assign MEM[34025] = MEM[806] + MEM[970];
assign MEM[34026] = MEM[810] + MEM[1407];
assign MEM[34027] = MEM[816] + MEM[1108];
assign MEM[34028] = MEM[821] + MEM[868];
assign MEM[34029] = MEM[829] + MEM[941];
assign MEM[34030] = MEM[842] + MEM[997];
assign MEM[34031] = MEM[844] + MEM[1294];
assign MEM[34032] = MEM[853] + MEM[1081];
assign MEM[34033] = MEM[854] + MEM[871];
assign MEM[34034] = MEM[855] + MEM[973];
assign MEM[34035] = MEM[863] + MEM[866];
assign MEM[34036] = MEM[870] + MEM[1023];
assign MEM[34037] = MEM[886] + MEM[902];
assign MEM[34038] = MEM[887] + MEM[1106];
assign MEM[34039] = MEM[911] + MEM[1109];
assign MEM[34040] = MEM[915] + MEM[1094];
assign MEM[34041] = MEM[917] + MEM[925];
assign MEM[34042] = MEM[931] + MEM[1058];
assign MEM[34043] = MEM[932] + MEM[1135];
assign MEM[34044] = MEM[934] + MEM[991];
assign MEM[34045] = MEM[942] + MEM[1309];
assign MEM[34046] = MEM[946] + MEM[1173];
assign MEM[34047] = MEM[948] + MEM[1406];
assign MEM[34048] = MEM[954] + MEM[1053];
assign MEM[34049] = MEM[956] + MEM[1034];
assign MEM[34050] = MEM[957] + MEM[1358];
assign MEM[34051] = MEM[958] + MEM[959];
assign MEM[34052] = MEM[960] + MEM[983];
assign MEM[34053] = MEM[964] + MEM[1671];
assign MEM[34054] = MEM[974] + MEM[1054];
assign MEM[34055] = MEM[986] + MEM[1044];
assign MEM[34056] = MEM[990] + MEM[1042];
assign MEM[34057] = MEM[994] + MEM[1455];
assign MEM[34058] = MEM[996] + MEM[1461];
assign MEM[34059] = MEM[1000] + MEM[1414];
assign MEM[34060] = MEM[1008] + MEM[1125];
assign MEM[34061] = MEM[1010] + MEM[1063];
assign MEM[34062] = MEM[1015] + MEM[1061];
assign MEM[34063] = MEM[1020] + MEM[1533];
assign MEM[34064] = MEM[1036] + MEM[1230];
assign MEM[34065] = MEM[1045] + MEM[1170];
assign MEM[34066] = MEM[1052] + MEM[1524];
assign MEM[34067] = MEM[1060] + MEM[1062];
assign MEM[34068] = MEM[1067] + MEM[1074];
assign MEM[34069] = MEM[1068] + MEM[1412];
assign MEM[34070] = MEM[1070] + MEM[1078];
assign MEM[34071] = MEM[1082] + MEM[1557];
assign MEM[34072] = MEM[1087] + MEM[1146];
assign MEM[34073] = MEM[1092] + MEM[1277];
assign MEM[34074] = MEM[1095] + MEM[1186];
assign MEM[34075] = MEM[1099] + MEM[1646];
assign MEM[34076] = MEM[1100] + MEM[1626];
assign MEM[34077] = MEM[1101] + MEM[1221];
assign MEM[34078] = MEM[1102] + MEM[1163];
assign MEM[34079] = MEM[1103] + MEM[1583];
assign MEM[34080] = MEM[1107] + MEM[1388];
assign MEM[34081] = MEM[1110] + MEM[1839];
assign MEM[34082] = MEM[1111] + MEM[1365];
assign MEM[34083] = MEM[1119] + MEM[1444];
assign MEM[34084] = MEM[1126] + MEM[1290];
assign MEM[34085] = MEM[1142] + MEM[1595];
assign MEM[34086] = MEM[1147] + MEM[1174];
assign MEM[34087] = MEM[1158] + MEM[1573];
assign MEM[34088] = MEM[1159] + MEM[1415];
assign MEM[34089] = MEM[1164] + MEM[1619];
assign MEM[34090] = MEM[1190] + MEM[1244];
assign MEM[34091] = MEM[1198] + MEM[1278];
assign MEM[34092] = MEM[1207] + MEM[1287];
assign MEM[34093] = MEM[1214] + MEM[1228];
assign MEM[34094] = MEM[1219] + MEM[1423];
assign MEM[34095] = MEM[1235] + MEM[1350];
assign MEM[34096] = MEM[1238] + MEM[1239];
assign MEM[34097] = MEM[1242] + MEM[1247];
assign MEM[34098] = MEM[1253] + MEM[1268];
assign MEM[34099] = MEM[1255] + MEM[1323];
assign MEM[34100] = MEM[1260] + MEM[1452];
assign MEM[34101] = MEM[1269] + MEM[1471];
assign MEM[34102] = MEM[1270] + MEM[1574];
assign MEM[34103] = MEM[1279] + MEM[1700];
assign MEM[34104] = MEM[1283] + MEM[1296];
assign MEM[34105] = MEM[1286] + MEM[1308];
assign MEM[34106] = MEM[1291] + MEM[1621];
assign MEM[34107] = MEM[1298] + MEM[1349];
assign MEM[34108] = MEM[1300] + MEM[1591];
assign MEM[34109] = MEM[1301] + MEM[1380];
assign MEM[34110] = MEM[1306] + MEM[1459];
assign MEM[34111] = MEM[1318] + MEM[1437];
assign MEM[34112] = MEM[1324] + MEM[1390];
assign MEM[34113] = MEM[1331] + MEM[1908];
assign MEM[34114] = MEM[1332] + MEM[1427];
assign MEM[34115] = MEM[1333] + MEM[1501];
assign MEM[34116] = MEM[1341] + MEM[1359];
assign MEM[34117] = MEM[1343] + MEM[1357];
assign MEM[34118] = MEM[1363] + MEM[1667];
assign MEM[34119] = MEM[1375] + MEM[1598];
assign MEM[34120] = MEM[1386] + MEM[1445];
assign MEM[34121] = MEM[1387] + MEM[2532];
assign MEM[34122] = MEM[1391] + MEM[1707];
assign MEM[34123] = MEM[1393] + MEM[2324];
assign MEM[34124] = MEM[1399] + MEM[1453];
assign MEM[34125] = MEM[1402] + MEM[1522];
assign MEM[34126] = MEM[1403] + MEM[1838];
assign MEM[34127] = MEM[1405] + MEM[1717];
assign MEM[34128] = MEM[1410] + MEM[1771];
assign MEM[34129] = MEM[1411] + MEM[1742];
assign MEM[34130] = MEM[1430] + MEM[1439];
assign MEM[34131] = MEM[1435] + MEM[1579];
assign MEM[34132] = MEM[1447] + MEM[1691];
assign MEM[34133] = MEM[1448] + MEM[1530];
assign MEM[34134] = MEM[1450] + MEM[1478];
assign MEM[34135] = MEM[1467] + MEM[1627];
assign MEM[34136] = MEM[1469] + MEM[1543];
assign MEM[34137] = MEM[1474] + MEM[1612];
assign MEM[34138] = MEM[1479] + MEM[1652];
assign MEM[34139] = MEM[1503] + MEM[1614];
assign MEM[34140] = MEM[1506] + MEM[1723];
assign MEM[34141] = MEM[1511] + MEM[1607];
assign MEM[34142] = MEM[1514] + MEM[1917];
assign MEM[34143] = MEM[1516] + MEM[1538];
assign MEM[34144] = MEM[1520] + MEM[1770];
assign MEM[34145] = MEM[1527] + MEM[1859];
assign MEM[34146] = MEM[1531] + MEM[1720];
assign MEM[34147] = MEM[1534] + MEM[1869];
assign MEM[34148] = MEM[1540] + MEM[1602];
assign MEM[34149] = MEM[1544] + MEM[1564];
assign MEM[34150] = MEM[1553] + MEM[1587];
assign MEM[34151] = MEM[1558] + MEM[2027];
assign MEM[34152] = MEM[1566] + MEM[1644];
assign MEM[34153] = MEM[1581] + MEM[1589];
assign MEM[34154] = MEM[1594] + MEM[1766];
assign MEM[34155] = MEM[1618] + MEM[1653];
assign MEM[34156] = MEM[1630] + MEM[1997];
assign MEM[34157] = MEM[1635] + MEM[1650];
assign MEM[34158] = MEM[1636] + MEM[1882];
assign MEM[34159] = MEM[1638] + MEM[1836];
assign MEM[34160] = MEM[1645] + MEM[1861];
assign MEM[34161] = MEM[1647] + MEM[1948];
assign MEM[34162] = MEM[1654] + MEM[1958];
assign MEM[34163] = MEM[1661] + MEM[1971];
assign MEM[34164] = MEM[1668] + MEM[1779];
assign MEM[34165] = MEM[1669] + MEM[1791];
assign MEM[34166] = MEM[1672] + MEM[1677];
assign MEM[34167] = MEM[1679] + MEM[1683];
assign MEM[34168] = MEM[1687] + MEM[1964];
assign MEM[34169] = MEM[1699] + MEM[1874];
assign MEM[34170] = MEM[1703] + MEM[1715];
assign MEM[34171] = MEM[1709] + MEM[1743];
assign MEM[34172] = MEM[1710] + MEM[3610];
assign MEM[34173] = MEM[1711] + MEM[2988];
assign MEM[34174] = MEM[1714] + MEM[2151];
assign MEM[34175] = MEM[1718] + MEM[1748];
assign MEM[34176] = MEM[1726] + MEM[1755];
assign MEM[34177] = MEM[1728] + MEM[1782];
assign MEM[34178] = MEM[1733] + MEM[1885];
assign MEM[34179] = MEM[1734] + MEM[2295];
assign MEM[34180] = MEM[1752] + MEM[1812];
assign MEM[34181] = MEM[1757] + MEM[1906];
assign MEM[34182] = MEM[1760] + MEM[1824];
assign MEM[34183] = MEM[1765] + MEM[2253];
assign MEM[34184] = MEM[1778] + MEM[1853];
assign MEM[34185] = MEM[1781] + MEM[2163];
assign MEM[34186] = MEM[1811] + MEM[2330];
assign MEM[34187] = MEM[1814] + MEM[1963];
assign MEM[34188] = MEM[1815] + MEM[2560];
assign MEM[34189] = MEM[1819] + MEM[2071];
assign MEM[34190] = MEM[1823] + MEM[1927];
assign MEM[34191] = MEM[1826] + MEM[1978];
assign MEM[34192] = MEM[1830] + MEM[1867];
assign MEM[34193] = MEM[1834] + MEM[1954];
assign MEM[34194] = MEM[1843] + MEM[2061];
assign MEM[34195] = MEM[1844] + MEM[2882];
assign MEM[34196] = MEM[1868] + MEM[1887];
assign MEM[34197] = MEM[1870] + MEM[1975];
assign MEM[34198] = MEM[1878] + MEM[2011];
assign MEM[34199] = MEM[1883] + MEM[2239];
assign MEM[34200] = MEM[1890] + MEM[2029];
assign MEM[34201] = MEM[1902] + MEM[2370];
assign MEM[34202] = MEM[1909] + MEM[1966];
assign MEM[34203] = MEM[1910] + MEM[1987];
assign MEM[34204] = MEM[1915] + MEM[2006];
assign MEM[34205] = MEM[1931] + MEM[1936];
assign MEM[34206] = MEM[1933] + MEM[1972];
assign MEM[34207] = MEM[1942] + MEM[2052];
assign MEM[34208] = MEM[1944] + MEM[1960];
assign MEM[34209] = MEM[1946] + MEM[2222];
assign MEM[34210] = MEM[1947] + MEM[2148];
assign MEM[34211] = MEM[1957] + MEM[2231];
assign MEM[34212] = MEM[1967] + MEM[2179];
assign MEM[34213] = MEM[1968] + MEM[2070];
assign MEM[34214] = MEM[1976] + MEM[2147];
assign MEM[34215] = MEM[1979] + MEM[2191];
assign MEM[34216] = MEM[1981] + MEM[2159];
assign MEM[34217] = MEM[1984] + MEM[2023];
assign MEM[34218] = MEM[1988] + MEM[2221];
assign MEM[34219] = MEM[1991] + MEM[2162];
assign MEM[34220] = MEM[1999] + MEM[2098];
assign MEM[34221] = MEM[2002] + MEM[2014];
assign MEM[34222] = MEM[2004] + MEM[2054];
assign MEM[34223] = MEM[2012] + MEM[2083];
assign MEM[34224] = MEM[2013] + MEM[2095];
assign MEM[34225] = MEM[2030] + MEM[2195];
assign MEM[34226] = MEM[2050] + MEM[2124];
assign MEM[34227] = MEM[2059] + MEM[2255];
assign MEM[34228] = MEM[2062] + MEM[2178];
assign MEM[34229] = MEM[2067] + MEM[2226];
assign MEM[34230] = MEM[2075] + MEM[2091];
assign MEM[34231] = MEM[2076] + MEM[2175];
assign MEM[34232] = MEM[2078] + MEM[2651];
assign MEM[34233] = MEM[2079] + MEM[2823];
assign MEM[34234] = MEM[2080] + MEM[2294];
assign MEM[34235] = MEM[2082] + MEM[2470];
assign MEM[34236] = MEM[2085] + MEM[2215];
assign MEM[34237] = MEM[2087] + MEM[2408];
assign MEM[34238] = MEM[2092] + MEM[2125];
assign MEM[34239] = MEM[2100] + MEM[2131];
assign MEM[34240] = MEM[2108] + MEM[2238];
assign MEM[34241] = MEM[2109] + MEM[2580];
assign MEM[34242] = MEM[2110] + MEM[2132];
assign MEM[34243] = MEM[2111] + MEM[2126];
assign MEM[34244] = MEM[2128] + MEM[2144];
assign MEM[34245] = MEM[2139] + MEM[2530];
assign MEM[34246] = MEM[2140] + MEM[2211];
assign MEM[34247] = MEM[2146] + MEM[2156];
assign MEM[34248] = MEM[2150] + MEM[2172];
assign MEM[34249] = MEM[2152] + MEM[2160];
assign MEM[34250] = MEM[2157] + MEM[2227];
assign MEM[34251] = MEM[2158] + MEM[2751];
assign MEM[34252] = MEM[2164] + MEM[2395];
assign MEM[34253] = MEM[2165] + MEM[2462];
assign MEM[34254] = MEM[2167] + MEM[2299];
assign MEM[34255] = MEM[2168] + MEM[2200];
assign MEM[34256] = MEM[2170] + MEM[2219];
assign MEM[34257] = MEM[2171] + MEM[2354];
assign MEM[34258] = MEM[2180] + MEM[2230];
assign MEM[34259] = MEM[2194] + MEM[2590];
assign MEM[34260] = MEM[2196] + MEM[2423];
assign MEM[34261] = MEM[2203] + MEM[2204];
assign MEM[34262] = MEM[2205] + MEM[2269];
assign MEM[34263] = MEM[2210] + MEM[2271];
assign MEM[34264] = MEM[2212] + MEM[2607];
assign MEM[34265] = MEM[2213] + MEM[2332];
assign MEM[34266] = MEM[2237] + MEM[2398];
assign MEM[34267] = MEM[2246] + MEM[2352];
assign MEM[34268] = MEM[2261] + MEM[2320];
assign MEM[34269] = MEM[2275] + MEM[2365];
assign MEM[34270] = MEM[2276] + MEM[2338];
assign MEM[34271] = MEM[2278] + MEM[2279];
assign MEM[34272] = MEM[2282] + MEM[2380];
assign MEM[34273] = MEM[2293] + MEM[2565];
assign MEM[34274] = MEM[2304] + MEM[2335];
assign MEM[34275] = MEM[2309] + MEM[2388];
assign MEM[34276] = MEM[2316] + MEM[2436];
assign MEM[34277] = MEM[2319] + MEM[2355];
assign MEM[34278] = MEM[2323] + MEM[2479];
assign MEM[34279] = MEM[2326] + MEM[2442];
assign MEM[34280] = MEM[2328] + MEM[2336];
assign MEM[34281] = MEM[2333] + MEM[2402];
assign MEM[34282] = MEM[2344] + MEM[2421];
assign MEM[34283] = MEM[2348] + MEM[2679];
assign MEM[34284] = MEM[2351] + MEM[2790];
assign MEM[34285] = MEM[2358] + MEM[2803];
assign MEM[34286] = MEM[2362] + MEM[2615];
assign MEM[34287] = MEM[2364] + MEM[2501];
assign MEM[34288] = MEM[2366] + MEM[2678];
assign MEM[34289] = MEM[2372] + MEM[2645];
assign MEM[34290] = MEM[2376] + MEM[2384];
assign MEM[34291] = MEM[2383] + MEM[2586];
assign MEM[34292] = MEM[2392] + MEM[2400];
assign MEM[34293] = MEM[2394] + MEM[2434];
assign MEM[34294] = MEM[2397] + MEM[2724];
assign MEM[34295] = MEM[2403] + MEM[2469];
assign MEM[34296] = MEM[2404] + MEM[2950];
assign MEM[34297] = MEM[2405] + MEM[2525];
assign MEM[34298] = MEM[2411] + MEM[2884];
assign MEM[34299] = MEM[2413] + MEM[2509];
assign MEM[34300] = MEM[2414] + MEM[2559];
assign MEM[34301] = MEM[2415] + MEM[3156];
assign MEM[34302] = MEM[2418] + MEM[2780];
assign MEM[34303] = MEM[2422] + MEM[2424];
assign MEM[34304] = MEM[2427] + MEM[2554];
assign MEM[34305] = MEM[2429] + MEM[2594];
assign MEM[34306] = MEM[2431] + MEM[2555];
assign MEM[34307] = MEM[2445] + MEM[2507];
assign MEM[34308] = MEM[2447] + MEM[2775];
assign MEM[34309] = MEM[2460] + MEM[2475];
assign MEM[34310] = MEM[2471] + MEM[3008];
assign MEM[34311] = MEM[2482] + MEM[2694];
assign MEM[34312] = MEM[2485] + MEM[2686];
assign MEM[34313] = MEM[2491] + MEM[2499];
assign MEM[34314] = MEM[2493] + MEM[2558];
assign MEM[34315] = MEM[2494] + MEM[2566];
assign MEM[34316] = MEM[2503] + MEM[2584];
assign MEM[34317] = MEM[2508] + MEM[2741];
assign MEM[34318] = MEM[2511] + MEM[2618];
assign MEM[34319] = MEM[2517] + MEM[2540];
assign MEM[34320] = MEM[2520] + MEM[2528];
assign MEM[34321] = MEM[2524] + MEM[2541];
assign MEM[34322] = MEM[2536] + MEM[2544];
assign MEM[34323] = MEM[2539] + MEM[2735];
assign MEM[34324] = MEM[2567] + MEM[2627];
assign MEM[34325] = MEM[2571] + MEM[2820];
assign MEM[34326] = MEM[2573] + MEM[2668];
assign MEM[34327] = MEM[2583] + MEM[3142];
assign MEM[34328] = MEM[2588] + MEM[2647];
assign MEM[34329] = MEM[2595] + MEM[2852];
assign MEM[34330] = MEM[2598] + MEM[2962];
assign MEM[34331] = MEM[2599] + MEM[2692];
assign MEM[34332] = MEM[2606] + MEM[2652];
assign MEM[34333] = MEM[2613] + MEM[2664];
assign MEM[34334] = MEM[2614] + MEM[2702];
assign MEM[34335] = MEM[2616] + MEM[2624];
assign MEM[34336] = MEM[2620] + MEM[2766];
assign MEM[34337] = MEM[2623] + MEM[2638];
assign MEM[34338] = MEM[2628] + MEM[2671];
assign MEM[34339] = MEM[2629] + MEM[2684];
assign MEM[34340] = MEM[2632] + MEM[2640];
assign MEM[34341] = MEM[2637] + MEM[2804];
assign MEM[34342] = MEM[2659] + MEM[2814];
assign MEM[34343] = MEM[2660] + MEM[2733];
assign MEM[34344] = MEM[2666] + MEM[2759];
assign MEM[34345] = MEM[2676] + MEM[2886];
assign MEM[34346] = MEM[2677] + MEM[2750];
assign MEM[34347] = MEM[2683] + MEM[2774];
assign MEM[34348] = MEM[2685] + MEM[3165];
assign MEM[34349] = MEM[2687] + MEM[2717];
assign MEM[34350] = MEM[2693] + MEM[2867];
assign MEM[34351] = MEM[2695] + MEM[3191];
assign MEM[34352] = MEM[2699] + MEM[2807];
assign MEM[34353] = MEM[2706] + MEM[2887];
assign MEM[34354] = MEM[2708] + MEM[2710];
assign MEM[34355] = MEM[2714] + MEM[2970];
assign MEM[34356] = MEM[2715] + MEM[2850];
assign MEM[34357] = MEM[2718] + MEM[2837];
assign MEM[34358] = MEM[2728] + MEM[2736];
assign MEM[34359] = MEM[2732] + MEM[2765];
assign MEM[34360] = MEM[2734] + MEM[2757];
assign MEM[34361] = MEM[2740] + MEM[2834];
assign MEM[34362] = MEM[2742] + MEM[2779];
assign MEM[34363] = MEM[2754] + MEM[3346];
assign MEM[34364] = MEM[2755] + MEM[3101];
assign MEM[34365] = MEM[2756] + MEM[2847];
assign MEM[34366] = MEM[2760] + MEM[2763];
assign MEM[34367] = MEM[2768] + MEM[2784];
assign MEM[34368] = MEM[2773] + MEM[3006];
assign MEM[34369] = MEM[2781] + MEM[2899];
assign MEM[34370] = MEM[2788] + MEM[3286];
assign MEM[34371] = MEM[2789] + MEM[2811];
assign MEM[34372] = MEM[2792] + MEM[2923];
assign MEM[34373] = MEM[2799] + MEM[2818];
assign MEM[34374] = MEM[2800] + MEM[2908];
assign MEM[34375] = MEM[2802] + MEM[2877];
assign MEM[34376] = MEM[2808] + MEM[2810];
assign MEM[34377] = MEM[2812] + MEM[2864];
assign MEM[34378] = MEM[2815] + MEM[2839];
assign MEM[34379] = MEM[2821] + MEM[2875];
assign MEM[34380] = MEM[2822] + MEM[3487];
assign MEM[34381] = MEM[2828] + MEM[2926];
assign MEM[34382] = MEM[2844] + MEM[3043];
assign MEM[34383] = MEM[2846] + MEM[2903];
assign MEM[34384] = MEM[2855] + MEM[3408];
assign MEM[34385] = MEM[2856] + MEM[2872];
assign MEM[34386] = MEM[2858] + MEM[3182];
assign MEM[34387] = MEM[2860] + MEM[2931];
assign MEM[34388] = MEM[2861] + MEM[3159];
assign MEM[34389] = MEM[2863] + MEM[2924];
assign MEM[34390] = MEM[2868] + MEM[3027];
assign MEM[34391] = MEM[2871] + MEM[2934];
assign MEM[34392] = MEM[2879] + MEM[3100];
assign MEM[34393] = MEM[2883] + MEM[2965];
assign MEM[34394] = MEM[2893] + MEM[2911];
assign MEM[34395] = MEM[2894] + MEM[2895];
assign MEM[34396] = MEM[2927] + MEM[2983];
assign MEM[34397] = MEM[2930] + MEM[3117];
assign MEM[34398] = MEM[2933] + MEM[2941];
assign MEM[34399] = MEM[2935] + MEM[3052];
assign MEM[34400] = MEM[2943] + MEM[2975];
assign MEM[34401] = MEM[2944] + MEM[2984];
assign MEM[34402] = MEM[2946] + MEM[3095];
assign MEM[34403] = MEM[2951] + MEM[3114];
assign MEM[34404] = MEM[2952] + MEM[3175];
assign MEM[34405] = MEM[2955] + MEM[3005];
assign MEM[34406] = MEM[2986] + MEM[3021];
assign MEM[34407] = MEM[2989] + MEM[3242];
assign MEM[34408] = MEM[2990] + MEM[3091];
assign MEM[34409] = MEM[2991] + MEM[3038];
assign MEM[34410] = MEM[2996] + MEM[3501];
assign MEM[34411] = MEM[2999] + MEM[3104];
assign MEM[34412] = MEM[3003] + MEM[3029];
assign MEM[34413] = MEM[3013] + MEM[3034];
assign MEM[34414] = MEM[3016] + MEM[3039];
assign MEM[34415] = MEM[3030] + MEM[3111];
assign MEM[34416] = MEM[3032] + MEM[3040];
assign MEM[34417] = MEM[3035] + MEM[3379];
assign MEM[34418] = MEM[3036] + MEM[3231];
assign MEM[34419] = MEM[3037] + MEM[3578];
assign MEM[34420] = MEM[3044] + MEM[3276];
assign MEM[34421] = MEM[3046] + MEM[3197];
assign MEM[34422] = MEM[3047] + MEM[3071];
assign MEM[34423] = MEM[3055] + MEM[3467];
assign MEM[34424] = MEM[3059] + MEM[3116];
assign MEM[34425] = MEM[3062] + MEM[3168];
assign MEM[34426] = MEM[3069] + MEM[3109];
assign MEM[34427] = MEM[3075] + MEM[3210];
assign MEM[34428] = MEM[3076] + MEM[3507];
assign MEM[34429] = MEM[3079] + MEM[3691];
assign MEM[34430] = MEM[3082] + MEM[3339];
assign MEM[34431] = MEM[3088] + MEM[3103];
assign MEM[34432] = MEM[3092] + MEM[3123];
assign MEM[34433] = MEM[3094] + MEM[3179];
assign MEM[34434] = MEM[3096] + MEM[3212];
assign MEM[34435] = MEM[3097] + MEM[3259];
assign MEM[34436] = MEM[3106] + MEM[3723];
assign MEM[34437] = MEM[3115] + MEM[3331];
assign MEM[34438] = MEM[3119] + MEM[3134];
assign MEM[34439] = MEM[3125] + MEM[3200];
assign MEM[34440] = MEM[3132] + MEM[3307];
assign MEM[34441] = MEM[3157] + MEM[4096];
assign MEM[34442] = MEM[3162] + MEM[3192];
assign MEM[34443] = MEM[3163] + MEM[3180];
assign MEM[34444] = MEM[3164] + MEM[3401];
assign MEM[34445] = MEM[3167] + MEM[3399];
assign MEM[34446] = MEM[3170] + MEM[3911];
assign MEM[34447] = MEM[3171] + MEM[3299];
assign MEM[34448] = MEM[3176] + MEM[3202];
assign MEM[34449] = MEM[3194] + MEM[3845];
assign MEM[34450] = MEM[3196] + MEM[3227];
assign MEM[34451] = MEM[3199] + MEM[3663];
assign MEM[34452] = MEM[3203] + MEM[3340];
assign MEM[34453] = MEM[3204] + MEM[3622];
assign MEM[34454] = MEM[3205] + MEM[3386];
assign MEM[34455] = MEM[3206] + MEM[3372];
assign MEM[34456] = MEM[3214] + MEM[3629];
assign MEM[34457] = MEM[3218] + MEM[3274];
assign MEM[34458] = MEM[3223] + MEM[3444];
assign MEM[34459] = MEM[3244] + MEM[3291];
assign MEM[34460] = MEM[3246] + MEM[3324];
assign MEM[34461] = MEM[3247] + MEM[3371];
assign MEM[34462] = MEM[3260] + MEM[3437];
assign MEM[34463] = MEM[3262] + MEM[3347];
assign MEM[34464] = MEM[3268] + MEM[3463];
assign MEM[34465] = MEM[3270] + MEM[3495];
assign MEM[34466] = MEM[3277] + MEM[3310];
assign MEM[34467] = MEM[3279] + MEM[3330];
assign MEM[34468] = MEM[3298] + MEM[3515];
assign MEM[34469] = MEM[3300] + MEM[3325];
assign MEM[34470] = MEM[3302] + MEM[3337];
assign MEM[34471] = MEM[3303] + MEM[3605];
assign MEM[34472] = MEM[3317] + MEM[3323];
assign MEM[34473] = MEM[3320] + MEM[3332];
assign MEM[34474] = MEM[3327] + MEM[3459];
assign MEM[34475] = MEM[3333] + MEM[3523];
assign MEM[34476] = MEM[3338] + MEM[3398];
assign MEM[34477] = MEM[3342] + MEM[3403];
assign MEM[34478] = MEM[3350] + MEM[3380];
assign MEM[34479] = MEM[3367] + MEM[3452];
assign MEM[34480] = MEM[3370] + MEM[3424];
assign MEM[34481] = MEM[3381] + MEM[3477];
assign MEM[34482] = MEM[3382] + MEM[3413];
assign MEM[34483] = MEM[3387] + MEM[3722];
assign MEM[34484] = MEM[3388] + MEM[3466];
assign MEM[34485] = MEM[3394] + MEM[3486];
assign MEM[34486] = MEM[3397] + MEM[3765];
assign MEM[34487] = MEM[3404] + MEM[3607];
assign MEM[34488] = MEM[3405] + MEM[4037];
assign MEM[34489] = MEM[3406] + MEM[3427];
assign MEM[34490] = MEM[3415] + MEM[3447];
assign MEM[34491] = MEM[3416] + MEM[3864];
assign MEM[34492] = MEM[3421] + MEM[3446];
assign MEM[34493] = MEM[3428] + MEM[3518];
assign MEM[34494] = MEM[3432] + MEM[3440];
assign MEM[34495] = MEM[3435] + MEM[3955];
assign MEM[34496] = MEM[3451] + MEM[3470];
assign MEM[34497] = MEM[3453] + MEM[3494];
assign MEM[34498] = MEM[3458] + MEM[3563];
assign MEM[34499] = MEM[3469] + MEM[3476];
assign MEM[34500] = MEM[3475] + MEM[3885];
assign MEM[34501] = MEM[3478] + MEM[3971];
assign MEM[34502] = MEM[3499] + MEM[3999];
assign MEM[34503] = MEM[3500] + MEM[3519];
assign MEM[34504] = MEM[3502] + MEM[3693];
assign MEM[34505] = MEM[3503] + MEM[3535];
assign MEM[34506] = MEM[3509] + MEM[3671];
assign MEM[34507] = MEM[3517] + MEM[3814];
assign MEM[34508] = MEM[3525] + MEM[3639];
assign MEM[34509] = MEM[3532] + MEM[3570];
assign MEM[34510] = MEM[3533] + MEM[3566];
assign MEM[34511] = MEM[3534] + MEM[3837];
assign MEM[34512] = MEM[3539] + MEM[3706];
assign MEM[34513] = MEM[3540] + MEM[3730];
assign MEM[34514] = MEM[3542] + MEM[3804];
assign MEM[34515] = MEM[3546] + MEM[3951];
assign MEM[34516] = MEM[3547] + MEM[4020];
assign MEM[34517] = MEM[3550] + MEM[3613];
assign MEM[34518] = MEM[3554] + MEM[3788];
assign MEM[34519] = MEM[3573] + MEM[3695];
assign MEM[34520] = MEM[3583] + MEM[3634];
assign MEM[34521] = MEM[3598] + MEM[3859];
assign MEM[34522] = MEM[3602] + MEM[3604];
assign MEM[34523] = MEM[3603] + MEM[3717];
assign MEM[34524] = MEM[3619] + MEM[3989];
assign MEM[34525] = MEM[3621] + MEM[3785];
assign MEM[34526] = MEM[3627] + MEM[3635];
assign MEM[34527] = MEM[3637] + MEM[3829];
assign MEM[34528] = MEM[3638] + MEM[3741];
assign MEM[34529] = MEM[3642] + MEM[3781];
assign MEM[34530] = MEM[3646] + MEM[3718];
assign MEM[34531] = MEM[3647] + MEM[3703];
assign MEM[34532] = MEM[3654] + MEM[3868];
assign MEM[34533] = MEM[3658] + MEM[4170];
assign MEM[34534] = MEM[3659] + MEM[3758];
assign MEM[34535] = MEM[3660] + MEM[3726];
assign MEM[34536] = MEM[3667] + MEM[3670];
assign MEM[34537] = MEM[3669] + MEM[3756];
assign MEM[34538] = MEM[3676] + MEM[3863];
assign MEM[34539] = MEM[3677] + MEM[3906];
assign MEM[34540] = MEM[3678] + MEM[3770];
assign MEM[34541] = MEM[3680] + MEM[3734];
assign MEM[34542] = MEM[3682] + MEM[3875];
assign MEM[34543] = MEM[3683] + MEM[3805];
assign MEM[34544] = MEM[3685] + MEM[4198];
assign MEM[34545] = MEM[3686] + MEM[3731];
assign MEM[34546] = MEM[3690] + MEM[3975];
assign MEM[34547] = MEM[3702] + MEM[3830];
assign MEM[34548] = MEM[3709] + MEM[3981];
assign MEM[34549] = MEM[3710] + MEM[3828];
assign MEM[34550] = MEM[3719] + MEM[3948];
assign MEM[34551] = MEM[3738] + MEM[3925];
assign MEM[34552] = MEM[3740] + MEM[3771];
assign MEM[34553] = MEM[3742] + MEM[3827];
assign MEM[34554] = MEM[3746] + MEM[4342];
assign MEM[34555] = MEM[3748] + MEM[3783];
assign MEM[34556] = MEM[3757] + MEM[3841];
assign MEM[34557] = MEM[3762] + MEM[3793];
assign MEM[34558] = MEM[3772] + MEM[4116];
assign MEM[34559] = MEM[3774] + MEM[3890];
assign MEM[34560] = MEM[3775] + MEM[3778];
assign MEM[34561] = MEM[3787] + MEM[3923];
assign MEM[34562] = MEM[3790] + MEM[3966];
assign MEM[34563] = MEM[3791] + MEM[3909];
assign MEM[34564] = MEM[3802] + MEM[3853];
assign MEM[34565] = MEM[3807] + MEM[3914];
assign MEM[34566] = MEM[3822] + MEM[3886];
assign MEM[34567] = MEM[3823] + MEM[4067];
assign MEM[34568] = MEM[3836] + MEM[3850];
assign MEM[34569] = MEM[3839] + MEM[4066];
assign MEM[34570] = MEM[3856] + MEM[4051];
assign MEM[34571] = MEM[3858] + MEM[4354];
assign MEM[34572] = MEM[3867] + MEM[3910];
assign MEM[34573] = MEM[3871] + MEM[3879];
assign MEM[34574] = MEM[3874] + MEM[4117];
assign MEM[34575] = MEM[3882] + MEM[4835];
assign MEM[34576] = MEM[3887] + MEM[3972];
assign MEM[34577] = MEM[3892] + MEM[3900];
assign MEM[34578] = MEM[3893] + MEM[4021];
assign MEM[34579] = MEM[3898] + MEM[3902];
assign MEM[34580] = MEM[3916] + MEM[4110];
assign MEM[34581] = MEM[3917] + MEM[4104];
assign MEM[34582] = MEM[3941] + MEM[4023];
assign MEM[34583] = MEM[3942] + MEM[4250];
assign MEM[34584] = MEM[3956] + MEM[3978];
assign MEM[34585] = MEM[3958] + MEM[4739];
assign MEM[34586] = MEM[3970] + MEM[4316];
assign MEM[34587] = MEM[3976] + MEM[3979];
assign MEM[34588] = MEM[3983] + MEM[4005];
assign MEM[34589] = MEM[3986] + MEM[4063];
assign MEM[34590] = MEM[3995] + MEM[4118];
assign MEM[34591] = MEM[3996] + MEM[4279];
assign MEM[34592] = MEM[3997] + MEM[4102];
assign MEM[34593] = MEM[4002] + MEM[4011];
assign MEM[34594] = MEM[4003] + MEM[4039];
assign MEM[34595] = MEM[4006] + MEM[4018];
assign MEM[34596] = MEM[4013] + MEM[4206];
assign MEM[34597] = MEM[4014] + MEM[4171];
assign MEM[34598] = MEM[4015] + MEM[4330];
assign MEM[34599] = MEM[4019] + MEM[4084];
assign MEM[34600] = MEM[4022] + MEM[4075];
assign MEM[34601] = MEM[4030] + MEM[4454];
assign MEM[34602] = MEM[4031] + MEM[4327];
assign MEM[34603] = MEM[4038] + MEM[4576];
assign MEM[34604] = MEM[4044] + MEM[4052];
assign MEM[34605] = MEM[4045] + MEM[4123];
assign MEM[34606] = MEM[4047] + MEM[4263];
assign MEM[34607] = MEM[4054] + MEM[4095];
assign MEM[34608] = MEM[4055] + MEM[4082];
assign MEM[34609] = MEM[4058] + MEM[4132];
assign MEM[34610] = MEM[4074] + MEM[4239];
assign MEM[34611] = MEM[4076] + MEM[4227];
assign MEM[34612] = MEM[4077] + MEM[4086];
assign MEM[34613] = MEM[4079] + MEM[4415];
assign MEM[34614] = MEM[4083] + MEM[4139];
assign MEM[34615] = MEM[4085] + MEM[4151];
assign MEM[34616] = MEM[4087] + MEM[4094];
assign MEM[34617] = MEM[4099] + MEM[4182];
assign MEM[34618] = MEM[4100] + MEM[4164];
assign MEM[34619] = MEM[4107] + MEM[4723];
assign MEM[34620] = MEM[4108] + MEM[4431];
assign MEM[34621] = MEM[4109] + MEM[4112];
assign MEM[34622] = MEM[4115] + MEM[4236];
assign MEM[34623] = MEM[4119] + MEM[4333];
assign MEM[34624] = MEM[4120] + MEM[4140];
assign MEM[34625] = MEM[4122] + MEM[4131];
assign MEM[34626] = MEM[4130] + MEM[4167];
assign MEM[34627] = MEM[4135] + MEM[4419];
assign MEM[34628] = MEM[4142] + MEM[4455];
assign MEM[34629] = MEM[4149] + MEM[4555];
assign MEM[34630] = MEM[4158] + MEM[4382];
assign MEM[34631] = MEM[4159] + MEM[4268];
assign MEM[34632] = MEM[4166] + MEM[4231];
assign MEM[34633] = MEM[4173] + MEM[4301];
assign MEM[34634] = MEM[4179] + MEM[4252];
assign MEM[34635] = MEM[4186] + MEM[4211];
assign MEM[34636] = MEM[4187] + MEM[4202];
assign MEM[34637] = MEM[4190] + MEM[4194];
assign MEM[34638] = MEM[4192] + MEM[4244];
assign MEM[34639] = MEM[4195] + MEM[4396];
assign MEM[34640] = MEM[4196] + MEM[4245];
assign MEM[34641] = MEM[4203] + MEM[4306];
assign MEM[34642] = MEM[4204] + MEM[4283];
assign MEM[34643] = MEM[4207] + MEM[4374];
assign MEM[34644] = MEM[4212] + MEM[4381];
assign MEM[34645] = MEM[4219] + MEM[4386];
assign MEM[34646] = MEM[4222] + MEM[4311];
assign MEM[34647] = MEM[4233] + MEM[4284];
assign MEM[34648] = MEM[4237] + MEM[4293];
assign MEM[34649] = MEM[4238] + MEM[4298];
assign MEM[34650] = MEM[4242] + MEM[4247];
assign MEM[34651] = MEM[4253] + MEM[4532];
assign MEM[34652] = MEM[4255] + MEM[4406];
assign MEM[34653] = MEM[4261] + MEM[4436];
assign MEM[34654] = MEM[4270] + MEM[4530];
assign MEM[34655] = MEM[4274] + MEM[4277];
assign MEM[34656] = MEM[4281] + MEM[4302];
assign MEM[34657] = MEM[4282] + MEM[4989];
assign MEM[34658] = MEM[4290] + MEM[4379];
assign MEM[34659] = MEM[4294] + MEM[4692];
assign MEM[34660] = MEM[4299] + MEM[4446];
assign MEM[34661] = MEM[4300] + MEM[4518];
assign MEM[34662] = MEM[4307] + MEM[4591];
assign MEM[34663] = MEM[4308] + MEM[4556];
assign MEM[34664] = MEM[4317] + MEM[4643];
assign MEM[34665] = MEM[4323] + MEM[4546];
assign MEM[34666] = MEM[4325] + MEM[4346];
assign MEM[34667] = MEM[4326] + MEM[4730];
assign MEM[34668] = MEM[4332] + MEM[4339];
assign MEM[34669] = MEM[4334] + MEM[4403];
assign MEM[34670] = MEM[4340] + MEM[4405];
assign MEM[34671] = MEM[4341] + MEM[4423];
assign MEM[34672] = MEM[4347] + MEM[4348];
assign MEM[34673] = MEM[4350] + MEM[4408];
assign MEM[34674] = MEM[4366] + MEM[4443];
assign MEM[34675] = MEM[4367] + MEM[4586];
assign MEM[34676] = MEM[4371] + MEM[4467];
assign MEM[34677] = MEM[4388] + MEM[4503];
assign MEM[34678] = MEM[4391] + MEM[4450];
assign MEM[34679] = MEM[4398] + MEM[5186];
assign MEM[34680] = MEM[4413] + MEM[4459];
assign MEM[34681] = MEM[4414] + MEM[4476];
assign MEM[34682] = MEM[4416] + MEM[4486];
assign MEM[34683] = MEM[4418] + MEM[4429];
assign MEM[34684] = MEM[4421] + MEM[4668];
assign MEM[34685] = MEM[4428] + MEM[4741];
assign MEM[34686] = MEM[4430] + MEM[5550];
assign MEM[34687] = MEM[4437] + MEM[4653];
assign MEM[34688] = MEM[4444] + MEM[4717];
assign MEM[34689] = MEM[4451] + MEM[4506];
assign MEM[34690] = MEM[4462] + MEM[4695];
assign MEM[34691] = MEM[4463] + MEM[4515];
assign MEM[34692] = MEM[4477] + MEM[4485];
assign MEM[34693] = MEM[4478] + MEM[5139];
assign MEM[34694] = MEM[4491] + MEM[4703];
assign MEM[34695] = MEM[4492] + MEM[4510];
assign MEM[34696] = MEM[4499] + MEM[4588];
assign MEM[34697] = MEM[4501] + MEM[4786];
assign MEM[34698] = MEM[4502] + MEM[4615];
assign MEM[34699] = MEM[4519] + MEM[4853];
assign MEM[34700] = MEM[4523] + MEM[4702];
assign MEM[34701] = MEM[4526] + MEM[4781];
assign MEM[34702] = MEM[4528] + MEM[4549];
assign MEM[34703] = MEM[4534] + MEM[4603];
assign MEM[34704] = MEM[4539] + MEM[4557];
assign MEM[34705] = MEM[4540] + MEM[5123];
assign MEM[34706] = MEM[4541] + MEM[5126];
assign MEM[34707] = MEM[4551] + MEM[4901];
assign MEM[34708] = MEM[4562] + MEM[4575];
assign MEM[34709] = MEM[4579] + MEM[4598];
assign MEM[34710] = MEM[4590] + MEM[4677];
assign MEM[34711] = MEM[4599] + MEM[4731];
assign MEM[34712] = MEM[4604] + MEM[4810];
assign MEM[34713] = MEM[4606] + MEM[4675];
assign MEM[34714] = MEM[4611] + MEM[4628];
assign MEM[34715] = MEM[4612] + MEM[4754];
assign MEM[34716] = MEM[4613] + MEM[4632];
assign MEM[34717] = MEM[4614] + MEM[4958];
assign MEM[34718] = MEM[4621] + MEM[4798];
assign MEM[34719] = MEM[4622] + MEM[5063];
assign MEM[34720] = MEM[4626] + MEM[4660];
assign MEM[34721] = MEM[4627] + MEM[4684];
assign MEM[34722] = MEM[4629] + MEM[4686];
assign MEM[34723] = MEM[4640] + MEM[4661];
assign MEM[34724] = MEM[4644] + MEM[4687];
assign MEM[34725] = MEM[4645] + MEM[4654];
assign MEM[34726] = MEM[4647] + MEM[4734];
assign MEM[34727] = MEM[4652] + MEM[4870];
assign MEM[34728] = MEM[4662] + MEM[4670];
assign MEM[34729] = MEM[4667] + MEM[4674];
assign MEM[34730] = MEM[4679] + MEM[4830];
assign MEM[34731] = MEM[4691] + MEM[5103];
assign MEM[34732] = MEM[4701] + MEM[5715];
assign MEM[34733] = MEM[4709] + MEM[4815];
assign MEM[34734] = MEM[4710] + MEM[4783];
assign MEM[34735] = MEM[4715] + MEM[4812];
assign MEM[34736] = MEM[4716] + MEM[5015];
assign MEM[34737] = MEM[4719] + MEM[4903];
assign MEM[34738] = MEM[4724] + MEM[5187];
assign MEM[34739] = MEM[4725] + MEM[5059];
assign MEM[34740] = MEM[4727] + MEM[4736];
assign MEM[34741] = MEM[4732] + MEM[6327];
assign MEM[34742] = MEM[4738] + MEM[4790];
assign MEM[34743] = MEM[4748] + MEM[4839];
assign MEM[34744] = MEM[4751] + MEM[4837];
assign MEM[34745] = MEM[4755] + MEM[4765];
assign MEM[34746] = MEM[4756] + MEM[5055];
assign MEM[34747] = MEM[4757] + MEM[4770];
assign MEM[34748] = MEM[4766] + MEM[5213];
assign MEM[34749] = MEM[4773] + MEM[4962];
assign MEM[34750] = MEM[4775] + MEM[4878];
assign MEM[34751] = MEM[4779] + MEM[4908];
assign MEM[34752] = MEM[4787] + MEM[4863];
assign MEM[34753] = MEM[4788] + MEM[4965];
assign MEM[34754] = MEM[4797] + MEM[4843];
assign MEM[34755] = MEM[4799] + MEM[4910];
assign MEM[34756] = MEM[4804] + MEM[4891];
assign MEM[34757] = MEM[4806] + MEM[5060];
assign MEM[34758] = MEM[4807] + MEM[4821];
assign MEM[34759] = MEM[4811] + MEM[4831];
assign MEM[34760] = MEM[4814] + MEM[5074];
assign MEM[34761] = MEM[4818] + MEM[4927];
assign MEM[34762] = MEM[4824] + MEM[5166];
assign MEM[34763] = MEM[4828] + MEM[5116];
assign MEM[34764] = MEM[4829] + MEM[4850];
assign MEM[34765] = MEM[4844] + MEM[4915];
assign MEM[34766] = MEM[4845] + MEM[4948];
assign MEM[34767] = MEM[4846] + MEM[4981];
assign MEM[34768] = MEM[4854] + MEM[4902];
assign MEM[34769] = MEM[4856] + MEM[5070];
assign MEM[34770] = MEM[4861] + MEM[5214];
assign MEM[34771] = MEM[4875] + MEM[4906];
assign MEM[34772] = MEM[4877] + MEM[5077];
assign MEM[34773] = MEM[4879] + MEM[4926];
assign MEM[34774] = MEM[4884] + MEM[4933];
assign MEM[34775] = MEM[4886] + MEM[4947];
assign MEM[34776] = MEM[4890] + MEM[5157];
assign MEM[34777] = MEM[4894] + MEM[5414];
assign MEM[34778] = MEM[4895] + MEM[5486];
assign MEM[34779] = MEM[4900] + MEM[5099];
assign MEM[34780] = MEM[4918] + MEM[4970];
assign MEM[34781] = MEM[4919] + MEM[4975];
assign MEM[34782] = MEM[4925] + MEM[4968];
assign MEM[34783] = MEM[4934] + MEM[5045];
assign MEM[34784] = MEM[4935] + MEM[5271];
assign MEM[34785] = MEM[4951] + MEM[5442];
assign MEM[34786] = MEM[4956] + MEM[4979];
assign MEM[34787] = MEM[4976] + MEM[4992];
assign MEM[34788] = MEM[4978] + MEM[5174];
assign MEM[34789] = MEM[4982] + MEM[5205];
assign MEM[34790] = MEM[4983] + MEM[5095];
assign MEM[34791] = MEM[4986] + MEM[5002];
assign MEM[34792] = MEM[4988] + MEM[5237];
assign MEM[34793] = MEM[4991] + MEM[5110];
assign MEM[34794] = MEM[4995] + MEM[5283];
assign MEM[34795] = MEM[4996] + MEM[5227];
assign MEM[34796] = MEM[4998] + MEM[5093];
assign MEM[34797] = MEM[4999] + MEM[5239];
assign MEM[34798] = MEM[5011] + MEM[5222];
assign MEM[34799] = MEM[5013] + MEM[5022];
assign MEM[34800] = MEM[5018] + MEM[5034];
assign MEM[34801] = MEM[5020] + MEM[5124];
assign MEM[34802] = MEM[5028] + MEM[5092];
assign MEM[34803] = MEM[5029] + MEM[5255];
assign MEM[34804] = MEM[5036] + MEM[5247];
assign MEM[34805] = MEM[5039] + MEM[5054];
assign MEM[34806] = MEM[5044] + MEM[5172];
assign MEM[34807] = MEM[5047] + MEM[5175];
assign MEM[34808] = MEM[5053] + MEM[5314];
assign MEM[34809] = MEM[5067] + MEM[5318];
assign MEM[34810] = MEM[5071] + MEM[5100];
assign MEM[34811] = MEM[5072] + MEM[5080];
assign MEM[34812] = MEM[5076] + MEM[5342];
assign MEM[34813] = MEM[5078] + MEM[5195];
assign MEM[34814] = MEM[5079] + MEM[5102];
assign MEM[34815] = MEM[5105] + MEM[5132];
assign MEM[34816] = MEM[5108] + MEM[5133];
assign MEM[34817] = MEM[5119] + MEM[5212];
assign MEM[34818] = MEM[5127] + MEM[5574];
assign MEM[34819] = MEM[5135] + MEM[5328];
assign MEM[34820] = MEM[5141] + MEM[5493];
assign MEM[34821] = MEM[5143] + MEM[5180];
assign MEM[34822] = MEM[5171] + MEM[5354];
assign MEM[34823] = MEM[5179] + MEM[5331];
assign MEM[34824] = MEM[5181] + MEM[5286];
assign MEM[34825] = MEM[5182] + MEM[5270];
assign MEM[34826] = MEM[5190] + MEM[5396];
assign MEM[34827] = MEM[5192] + MEM[5250];
assign MEM[34828] = MEM[5199] + MEM[5335];
assign MEM[34829] = MEM[5203] + MEM[5432];
assign MEM[34830] = MEM[5204] + MEM[5333];
assign MEM[34831] = MEM[5229] + MEM[5629];
assign MEM[34832] = MEM[5230] + MEM[5412];
assign MEM[34833] = MEM[5234] + MEM[5242];
assign MEM[34834] = MEM[5243] + MEM[5346];
assign MEM[34835] = MEM[5244] + MEM[5750];
assign MEM[34836] = MEM[5252] + MEM[5435];
assign MEM[34837] = MEM[5261] + MEM[5307];
assign MEM[34838] = MEM[5263] + MEM[5781];
assign MEM[34839] = MEM[5277] + MEM[5296];
assign MEM[34840] = MEM[5278] + MEM[5397];
assign MEM[34841] = MEM[5279] + MEM[5572];
assign MEM[34842] = MEM[5280] + MEM[5496];
assign MEM[34843] = MEM[5287] + MEM[5695];
assign MEM[34844] = MEM[5290] + MEM[5846];
assign MEM[34845] = MEM[5291] + MEM[5340];
assign MEM[34846] = MEM[5292] + MEM[5487];
assign MEM[34847] = MEM[5295] + MEM[5437];
assign MEM[34848] = MEM[5303] + MEM[5419];
assign MEM[34849] = MEM[5308] + MEM[5319];
assign MEM[34850] = MEM[5309] + MEM[5698];
assign MEM[34851] = MEM[5310] + MEM[5778];
assign MEM[34852] = MEM[5317] + MEM[5334];
assign MEM[34853] = MEM[5321] + MEM[5338];
assign MEM[34854] = MEM[5322] + MEM[5363];
assign MEM[34855] = MEM[5324] + MEM[5566];
assign MEM[34856] = MEM[5327] + MEM[5977];
assign MEM[34857] = MEM[5350] + MEM[5658];
assign MEM[34858] = MEM[5355] + MEM[5438];
assign MEM[34859] = MEM[5357] + MEM[5559];
assign MEM[34860] = MEM[5359] + MEM[5444];
assign MEM[34861] = MEM[5364] + MEM[5742];
assign MEM[34862] = MEM[5366] + MEM[5506];
assign MEM[34863] = MEM[5367] + MEM[5542];
assign MEM[34864] = MEM[5374] + MEM[5445];
assign MEM[34865] = MEM[5391] + MEM[5431];
assign MEM[34866] = MEM[5398] + MEM[5454];
assign MEM[34867] = MEM[5403] + MEM[5409];
assign MEM[34868] = MEM[5406] + MEM[5508];
assign MEM[34869] = MEM[5407] + MEM[5478];
assign MEM[34870] = MEM[5410] + MEM[5458];
assign MEM[34871] = MEM[5411] + MEM[5663];
assign MEM[34872] = MEM[5415] + MEM[5651];
assign MEM[34873] = MEM[5420] + MEM[5453];
assign MEM[34874] = MEM[5424] + MEM[5426];
assign MEM[34875] = MEM[5427] + MEM[5759];
assign MEM[34876] = MEM[5440] + MEM[5744];
assign MEM[34877] = MEM[5450] + MEM[5510];
assign MEM[34878] = MEM[5463] + MEM[5466];
assign MEM[34879] = MEM[5467] + MEM[5719];
assign MEM[34880] = MEM[5476] + MEM[5644];
assign MEM[34881] = MEM[5484] + MEM[5755];
assign MEM[34882] = MEM[5491] + MEM[5551];
assign MEM[34883] = MEM[5492] + MEM[5718];
assign MEM[34884] = MEM[5495] + MEM[5887];
assign MEM[34885] = MEM[5501] + MEM[5733];
assign MEM[34886] = MEM[5502] + MEM[5562];
assign MEM[34887] = MEM[5503] + MEM[5736];
assign MEM[34888] = MEM[5504] + MEM[5691];
assign MEM[34889] = MEM[5509] + MEM[5948];
assign MEM[34890] = MEM[5518] + MEM[5525];
assign MEM[34891] = MEM[5519] + MEM[5866];
assign MEM[34892] = MEM[5522] + MEM[5726];
assign MEM[34893] = MEM[5532] + MEM[5700];
assign MEM[34894] = MEM[5537] + MEM[5541];
assign MEM[34895] = MEM[5538] + MEM[5790];
assign MEM[34896] = MEM[5539] + MEM[5746];
assign MEM[34897] = MEM[5548] + MEM[5735];
assign MEM[34898] = MEM[5557] + MEM[6071];
assign MEM[34899] = MEM[5563] + MEM[5660];
assign MEM[34900] = MEM[5564] + MEM[5712];
assign MEM[34901] = MEM[5567] + MEM[5679];
assign MEM[34902] = MEM[5575] + MEM[5752];
assign MEM[34903] = MEM[5579] + MEM[5647];
assign MEM[34904] = MEM[5581] + MEM[5787];
assign MEM[34905] = MEM[5590] + MEM[5957];
assign MEM[34906] = MEM[5605] + MEM[5607];
assign MEM[34907] = MEM[5628] + MEM[5675];
assign MEM[34908] = MEM[5630] + MEM[5636];
assign MEM[34909] = MEM[5639] + MEM[5783];
assign MEM[34910] = MEM[5649] + MEM[5665];
assign MEM[34911] = MEM[5653] + MEM[5771];
assign MEM[34912] = MEM[5654] + MEM[5725];
assign MEM[34913] = MEM[5670] + MEM[5724];
assign MEM[34914] = MEM[5671] + MEM[5687];
assign MEM[34915] = MEM[5677] + MEM[6472];
assign MEM[34916] = MEM[5683] + MEM[5749];
assign MEM[34917] = MEM[5686] + MEM[5709];
assign MEM[34918] = MEM[5690] + MEM[5732];
assign MEM[34919] = MEM[5701] + MEM[5868];
assign MEM[34920] = MEM[5706] + MEM[5743];
assign MEM[34921] = MEM[5708] + MEM[5916];
assign MEM[34922] = MEM[5714] + MEM[5767];
assign MEM[34923] = MEM[5728] + MEM[5730];
assign MEM[34924] = MEM[5731] + MEM[5814];
assign MEM[34925] = MEM[5737] + MEM[5738];
assign MEM[34926] = MEM[5739] + MEM[5741];
assign MEM[34927] = MEM[5740] + MEM[6167];
assign MEM[34928] = MEM[5751] + MEM[6126];
assign MEM[34929] = MEM[5757] + MEM[5799];
assign MEM[34930] = MEM[5765] + MEM[5775];
assign MEM[34931] = MEM[5772] + MEM[5946];
assign MEM[34932] = MEM[5779] + MEM[5854];
assign MEM[34933] = MEM[5788] + MEM[5805];
assign MEM[34934] = MEM[5789] + MEM[6405];
assign MEM[34935] = MEM[5791] + MEM[5796];
assign MEM[34936] = MEM[5797] + MEM[5927];
assign MEM[34937] = MEM[5829] + MEM[5935];
assign MEM[34938] = MEM[5838] + MEM[6015];
assign MEM[34939] = MEM[5858] + MEM[5876];
assign MEM[34940] = MEM[5859] + MEM[5879];
assign MEM[34941] = MEM[5863] + MEM[5902];
assign MEM[34942] = MEM[5867] + MEM[6037];
assign MEM[34943] = MEM[5871] + MEM[6150];
assign MEM[34944] = MEM[5874] + MEM[6269];
assign MEM[34945] = MEM[5877] + MEM[5951];
assign MEM[34946] = MEM[5878] + MEM[5994];
assign MEM[34947] = MEM[5882] + MEM[6283];
assign MEM[34948] = MEM[5885] + MEM[5918];
assign MEM[34949] = MEM[5886] + MEM[5936];
assign MEM[34950] = MEM[5890] + MEM[6367];
assign MEM[34951] = MEM[5891] + MEM[5974];
assign MEM[34952] = MEM[5893] + MEM[6294];
assign MEM[34953] = MEM[5898] + MEM[5904];
assign MEM[34954] = MEM[5906] + MEM[6101];
assign MEM[34955] = MEM[5908] + MEM[5999];
assign MEM[34956] = MEM[5910] + MEM[5972];
assign MEM[34957] = MEM[5912] + MEM[6183];
assign MEM[34958] = MEM[5919] + MEM[6002];
assign MEM[34959] = MEM[5926] + MEM[5942];
assign MEM[34960] = MEM[5929] + MEM[6334];
assign MEM[34961] = MEM[5930] + MEM[6370];
assign MEM[34962] = MEM[5931] + MEM[5947];
assign MEM[34963] = MEM[5932] + MEM[5968];
assign MEM[34964] = MEM[5941] + MEM[5950];
assign MEM[34965] = MEM[5944] + MEM[6138];
assign MEM[34966] = MEM[5954] + MEM[6093];
assign MEM[34967] = MEM[5955] + MEM[6422];
assign MEM[34968] = MEM[5964] + MEM[6203];
assign MEM[34969] = MEM[5965] + MEM[6379];
assign MEM[34970] = MEM[5967] + MEM[5978];
assign MEM[34971] = MEM[5971] + MEM[6142];
assign MEM[34972] = MEM[5979] + MEM[6154];
assign MEM[34973] = MEM[5980] + MEM[6817];
assign MEM[34974] = MEM[5981] + MEM[6124];
assign MEM[34975] = MEM[5982] + MEM[6668];
assign MEM[34976] = MEM[5988] + MEM[6725];
assign MEM[34977] = MEM[5995] + MEM[6095];
assign MEM[34978] = MEM[5996] + MEM[6143];
assign MEM[34979] = MEM[5997] + MEM[6061];
assign MEM[34980] = MEM[5998] + MEM[6419];
assign MEM[34981] = MEM[6003] + MEM[6310];
assign MEM[34982] = MEM[6007] + MEM[6672];
assign MEM[34983] = MEM[6012] + MEM[6173];
assign MEM[34984] = MEM[6013] + MEM[6221];
assign MEM[34985] = MEM[6022] + MEM[6212];
assign MEM[34986] = MEM[6039] + MEM[6309];
assign MEM[34987] = MEM[6055] + MEM[6070];
assign MEM[34988] = MEM[6062] + MEM[6108];
assign MEM[34989] = MEM[6063] + MEM[6155];
assign MEM[34990] = MEM[6079] + MEM[6273];
assign MEM[34991] = MEM[6086] + MEM[6179];
assign MEM[34992] = MEM[6102] + MEM[6110];
assign MEM[34993] = MEM[6103] + MEM[6199];
assign MEM[34994] = MEM[6107] + MEM[6156];
assign MEM[34995] = MEM[6133] + MEM[6162];
assign MEM[34996] = MEM[6134] + MEM[6276];
assign MEM[34997] = MEM[6140] + MEM[6388];
assign MEM[34998] = MEM[6147] + MEM[6151];
assign MEM[34999] = MEM[6158] + MEM[6425];
assign MEM[35000] = MEM[6164] + MEM[6468];
assign MEM[35001] = MEM[6178] + MEM[6620];
assign MEM[35002] = MEM[6187] + MEM[6190];
assign MEM[35003] = MEM[6196] + MEM[6281];
assign MEM[35004] = MEM[6197] + MEM[6230];
assign MEM[35005] = MEM[6206] + MEM[6361];
assign MEM[35006] = MEM[6222] + MEM[6358];
assign MEM[35007] = MEM[6228] + MEM[6430];
assign MEM[35008] = MEM[6231] + MEM[6446];
assign MEM[35009] = MEM[6247] + MEM[6420];
assign MEM[35010] = MEM[6263] + MEM[6270];
assign MEM[35011] = MEM[6274] + MEM[6373];
assign MEM[35012] = MEM[6275] + MEM[6538];
assign MEM[35013] = MEM[6277] + MEM[6335];
assign MEM[35014] = MEM[6287] + MEM[6295];
assign MEM[35015] = MEM[6288] + MEM[6752];
assign MEM[35016] = MEM[6291] + MEM[6365];
assign MEM[35017] = MEM[6293] + MEM[6484];
assign MEM[35018] = MEM[6298] + MEM[6333];
assign MEM[35019] = MEM[6300] + MEM[6313];
assign MEM[35020] = MEM[6301] + MEM[6863];
assign MEM[35021] = MEM[6303] + MEM[6429];
assign MEM[35022] = MEM[6304] + MEM[6353];
assign MEM[35023] = MEM[6311] + MEM[6345];
assign MEM[35024] = MEM[6318] + MEM[6423];
assign MEM[35025] = MEM[6322] + MEM[7497];
assign MEM[35026] = MEM[6332] + MEM[6427];
assign MEM[35027] = MEM[6337] + MEM[6340];
assign MEM[35028] = MEM[6339] + MEM[6377];
assign MEM[35029] = MEM[6341] + MEM[6798];
assign MEM[35030] = MEM[6342] + MEM[6362];
assign MEM[35031] = MEM[6346] + MEM[6385];
assign MEM[35032] = MEM[6347] + MEM[6413];
assign MEM[35033] = MEM[6360] + MEM[6390];
assign MEM[35034] = MEM[6363] + MEM[6849];
assign MEM[35035] = MEM[6369] + MEM[6709];
assign MEM[35036] = MEM[6374] + MEM[6519];
assign MEM[35037] = MEM[6376] + MEM[6424];
assign MEM[35038] = MEM[6402] + MEM[6516];
assign MEM[35039] = MEM[6412] + MEM[6948];
assign MEM[35040] = MEM[6414] + MEM[6505];
assign MEM[35041] = MEM[6426] + MEM[6915];
assign MEM[35042] = MEM[6432] + MEM[6547];
assign MEM[35043] = MEM[6435] + MEM[6975];
assign MEM[35044] = MEM[6441] + MEM[6501];
assign MEM[35045] = MEM[6444] + MEM[6493];
assign MEM[35046] = MEM[6455] + MEM[6488];
assign MEM[35047] = MEM[6463] + MEM[6506];
assign MEM[35048] = MEM[6464] + MEM[6657];
assign MEM[35049] = MEM[6465] + MEM[6480];
assign MEM[35050] = MEM[6476] + MEM[6660];
assign MEM[35051] = MEM[6478] + MEM[6525];
assign MEM[35052] = MEM[6492] + MEM[6584];
assign MEM[35053] = MEM[6494] + MEM[6614];
assign MEM[35054] = MEM[6495] + MEM[6598];
assign MEM[35055] = MEM[6497] + MEM[6524];
assign MEM[35056] = MEM[6498] + MEM[6499];
assign MEM[35057] = MEM[6512] + MEM[6523];
assign MEM[35058] = MEM[6514] + MEM[6631];
assign MEM[35059] = MEM[6536] + MEM[6613];
assign MEM[35060] = MEM[6546] + MEM[6897];
assign MEM[35061] = MEM[6548] + MEM[6696];
assign MEM[35062] = MEM[6559] + MEM[6679];
assign MEM[35063] = MEM[6561] + MEM[6563];
assign MEM[35064] = MEM[6564] + MEM[6615];
assign MEM[35065] = MEM[6569] + MEM[6636];
assign MEM[35066] = MEM[6570] + MEM[6976];
assign MEM[35067] = MEM[6571] + MEM[6612];
assign MEM[35068] = MEM[6579] + MEM[6588];
assign MEM[35069] = MEM[6582] + MEM[6706];
assign MEM[35070] = MEM[6585] + MEM[6847];
assign MEM[35071] = MEM[6589] + MEM[6916];
assign MEM[35072] = MEM[6590] + MEM[7099];
assign MEM[35073] = MEM[6591] + MEM[6617];
assign MEM[35074] = MEM[6608] + MEM[6903];
assign MEM[35075] = MEM[6619] + MEM[6658];
assign MEM[35076] = MEM[6629] + MEM[6716];
assign MEM[35077] = MEM[6633] + MEM[6714];
assign MEM[35078] = MEM[6651] + MEM[6701];
assign MEM[35079] = MEM[6659] + MEM[6718];
assign MEM[35080] = MEM[6663] + MEM[6747];
assign MEM[35081] = MEM[6669] + MEM[6871];
assign MEM[35082] = MEM[6675] + MEM[6681];
assign MEM[35083] = MEM[6678] + MEM[6901];
assign MEM[35084] = MEM[6695] + MEM[6787];
assign MEM[35085] = MEM[6697] + MEM[7711];
assign MEM[35086] = MEM[6699] + MEM[6831];
assign MEM[35087] = MEM[6702] + MEM[6874];
assign MEM[35088] = MEM[6708] + MEM[6992];
assign MEM[35089] = MEM[6710] + MEM[6723];
assign MEM[35090] = MEM[6724] + MEM[7213];
assign MEM[35091] = MEM[6738] + MEM[6879];
assign MEM[35092] = MEM[6743] + MEM[6806];
assign MEM[35093] = MEM[6748] + MEM[6812];
assign MEM[35094] = MEM[6750] + MEM[6913];
assign MEM[35095] = MEM[6775] + MEM[7159];
assign MEM[35096] = MEM[6779] + MEM[7259];
assign MEM[35097] = MEM[6784] + MEM[6900];
assign MEM[35098] = MEM[6795] + MEM[6922];
assign MEM[35099] = MEM[6796] + MEM[6842];
assign MEM[35100] = MEM[6797] + MEM[6844];
assign MEM[35101] = MEM[6799] + MEM[7208];
assign MEM[35102] = MEM[6803] + MEM[7335];
assign MEM[35103] = MEM[6804] + MEM[6873];
assign MEM[35104] = MEM[6807] + MEM[7161];
assign MEM[35105] = MEM[6808] + MEM[7034];
assign MEM[35106] = MEM[6809] + MEM[6906];
assign MEM[35107] = MEM[6813] + MEM[7144];
assign MEM[35108] = MEM[6814] + MEM[6930];
assign MEM[35109] = MEM[6816] + MEM[7109];
assign MEM[35110] = MEM[6819] + MEM[6857];
assign MEM[35111] = MEM[6821] + MEM[6955];
assign MEM[35112] = MEM[6832] + MEM[7308];
assign MEM[35113] = MEM[6836] + MEM[6937];
assign MEM[35114] = MEM[6838] + MEM[6957];
assign MEM[35115] = MEM[6859] + MEM[6899];
assign MEM[35116] = MEM[6866] + MEM[7025];
assign MEM[35117] = MEM[6876] + MEM[6954];
assign MEM[35118] = MEM[6886] + MEM[6921];
assign MEM[35119] = MEM[6887] + MEM[6889];
assign MEM[35120] = MEM[6905] + MEM[7022];
assign MEM[35121] = MEM[6908] + MEM[7217];
assign MEM[35122] = MEM[6914] + MEM[7073];
assign MEM[35123] = MEM[6928] + MEM[6980];
assign MEM[35124] = MEM[6929] + MEM[7479];
assign MEM[35125] = MEM[6933] + MEM[7035];
assign MEM[35126] = MEM[6942] + MEM[7013];
assign MEM[35127] = MEM[6943] + MEM[7224];
assign MEM[35128] = MEM[6944] + MEM[7333];
assign MEM[35129] = MEM[6951] + MEM[7088];
assign MEM[35130] = MEM[6952] + MEM[7495];
assign MEM[35131] = MEM[6959] + MEM[7143];
assign MEM[35132] = MEM[6973] + MEM[7110];
assign MEM[35133] = MEM[6984] + MEM[7005];
assign MEM[35134] = MEM[6985] + MEM[7037];
assign MEM[35135] = MEM[6987] + MEM[7269];
assign MEM[35136] = MEM[6995] + MEM[6996];
assign MEM[35137] = MEM[7001] + MEM[7074];
assign MEM[35138] = MEM[7006] + MEM[7209];
assign MEM[35139] = MEM[7015] + MEM[7021];
assign MEM[35140] = MEM[7019] + MEM[7172];
assign MEM[35141] = MEM[7023] + MEM[7171];
assign MEM[35142] = MEM[7026] + MEM[7084];
assign MEM[35143] = MEM[7027] + MEM[7112];
assign MEM[35144] = MEM[7028] + MEM[7193];
assign MEM[35145] = MEM[7029] + MEM[7046];
assign MEM[35146] = MEM[7038] + MEM[7106];
assign MEM[35147] = MEM[7042] + MEM[7051];
assign MEM[35148] = MEM[7048] + MEM[7139];
assign MEM[35149] = MEM[7050] + MEM[7243];
assign MEM[35150] = MEM[7052] + MEM[7297];
assign MEM[35151] = MEM[7053] + MEM[7280];
assign MEM[35152] = MEM[7054] + MEM[7097];
assign MEM[35153] = MEM[7055] + MEM[7986];
assign MEM[35154] = MEM[7056] + MEM[7184];
assign MEM[35155] = MEM[7062] + MEM[7151];
assign MEM[35156] = MEM[7065] + MEM[7180];
assign MEM[35157] = MEM[7076] + MEM[7141];
assign MEM[35158] = MEM[7083] + MEM[7392];
assign MEM[35159] = MEM[7094] + MEM[7275];
assign MEM[35160] = MEM[7102] + MEM[7165];
assign MEM[35161] = MEM[7105] + MEM[7292];
assign MEM[35162] = MEM[7115] + MEM[7129];
assign MEM[35163] = MEM[7117] + MEM[7211];
assign MEM[35164] = MEM[7118] + MEM[7200];
assign MEM[35165] = MEM[7120] + MEM[7359];
assign MEM[35166] = MEM[7123] + MEM[7307];
assign MEM[35167] = MEM[7126] + MEM[7703];
assign MEM[35168] = MEM[7130] + MEM[7142];
assign MEM[35169] = MEM[7133] + MEM[7278];
assign MEM[35170] = MEM[7137] + MEM[7199];
assign MEM[35171] = MEM[7140] + MEM[7241];
assign MEM[35172] = MEM[7147] + MEM[7216];
assign MEM[35173] = MEM[7162] + MEM[7414];
assign MEM[35174] = MEM[7169] + MEM[7179];
assign MEM[35175] = MEM[7175] + MEM[7233];
assign MEM[35176] = MEM[7176] + MEM[7237];
assign MEM[35177] = MEM[7178] + MEM[7363];
assign MEM[35178] = MEM[7192] + MEM[7261];
assign MEM[35179] = MEM[7202] + MEM[7646];
assign MEM[35180] = MEM[7206] + MEM[7337];
assign MEM[35181] = MEM[7212] + MEM[7423];
assign MEM[35182] = MEM[7219] + MEM[7357];
assign MEM[35183] = MEM[7225] + MEM[7382];
assign MEM[35184] = MEM[7234] + MEM[7388];
assign MEM[35185] = MEM[7235] + MEM[7242];
assign MEM[35186] = MEM[7244] + MEM[7287];
assign MEM[35187] = MEM[7247] + MEM[7311];
assign MEM[35188] = MEM[7254] + MEM[7282];
assign MEM[35189] = MEM[7260] + MEM[7290];
assign MEM[35190] = MEM[7276] + MEM[7344];
assign MEM[35191] = MEM[7284] + MEM[7293];
assign MEM[35192] = MEM[7285] + MEM[7451];
assign MEM[35193] = MEM[7288] + MEM[7478];
assign MEM[35194] = MEM[7289] + MEM[7390];
assign MEM[35195] = MEM[7291] + MEM[7693];
assign MEM[35196] = MEM[7296] + MEM[7430];
assign MEM[35197] = MEM[7299] + MEM[7802];
assign MEM[35198] = MEM[7300] + MEM[7312];
assign MEM[35199] = MEM[7301] + MEM[7321];
assign MEM[35200] = MEM[7302] + MEM[7593];
assign MEM[35201] = MEM[7304] + MEM[7486];
assign MEM[35202] = MEM[7305] + MEM[7374];
assign MEM[35203] = MEM[7306] + MEM[7580];
assign MEM[35204] = MEM[7310] + MEM[7383];
assign MEM[35205] = MEM[7318] + MEM[7351];
assign MEM[35206] = MEM[7322] + MEM[7331];
assign MEM[35207] = MEM[7325] + MEM[7463];
assign MEM[35208] = MEM[7332] + MEM[7483];
assign MEM[35209] = MEM[7338] + MEM[7413];
assign MEM[35210] = MEM[7339] + MEM[7441];
assign MEM[35211] = MEM[7340] + MEM[7381];
assign MEM[35212] = MEM[7341] + MEM[7438];
assign MEM[35213] = MEM[7342] + MEM[7472];
assign MEM[35214] = MEM[7352] + MEM[7371];
assign MEM[35215] = MEM[7354] + MEM[7454];
assign MEM[35216] = MEM[7369] + MEM[7534];
assign MEM[35217] = MEM[7380] + MEM[7410];
assign MEM[35218] = MEM[7385] + MEM[7386];
assign MEM[35219] = MEM[7394] + MEM[7428];
assign MEM[35220] = MEM[7399] + MEM[7469];
assign MEM[35221] = MEM[7420] + MEM[7546];
assign MEM[35222] = MEM[7429] + MEM[7686];
assign MEM[35223] = MEM[7433] + MEM[7532];
assign MEM[35224] = MEM[7439] + MEM[7966];
assign MEM[35225] = MEM[7443] + MEM[7648];
assign MEM[35226] = MEM[7452] + MEM[7523];
assign MEM[35227] = MEM[7455] + MEM[7490];
assign MEM[35228] = MEM[7457] + MEM[7531];
assign MEM[35229] = MEM[7458] + MEM[7567];
assign MEM[35230] = MEM[7459] + MEM[7539];
assign MEM[35231] = MEM[7462] + MEM[7615];
assign MEM[35232] = MEM[7477] + MEM[7491];
assign MEM[35233] = MEM[7480] + MEM[7590];
assign MEM[35234] = MEM[7489] + MEM[7676];
assign MEM[35235] = MEM[7498] + MEM[7545];
assign MEM[35236] = MEM[7500] + MEM[7649];
assign MEM[35237] = MEM[7502] + MEM[7685];
assign MEM[35238] = MEM[7503] + MEM[7674];
assign MEM[35239] = MEM[7505] + MEM[7767];
assign MEM[35240] = MEM[7508] + MEM[7653];
assign MEM[35241] = MEM[7511] + MEM[7652];
assign MEM[35242] = MEM[7512] + MEM[7737];
assign MEM[35243] = MEM[7528] + MEM[7914];
assign MEM[35244] = MEM[7537] + MEM[7763];
assign MEM[35245] = MEM[7538] + MEM[7560];
assign MEM[35246] = MEM[7540] + MEM[7610];
assign MEM[35247] = MEM[7542] + MEM[7806];
assign MEM[35248] = MEM[7543] + MEM[7597];
assign MEM[35249] = MEM[7550] + MEM[7816];
assign MEM[35250] = MEM[7552] + MEM[7571];
assign MEM[35251] = MEM[7566] + MEM[7882];
assign MEM[35252] = MEM[7570] + MEM[7614];
assign MEM[35253] = MEM[7576] + MEM[7951];
assign MEM[35254] = MEM[7577] + MEM[7672];
assign MEM[35255] = MEM[7581] + MEM[7886];
assign MEM[35256] = MEM[7592] + MEM[7715];
assign MEM[35257] = MEM[7594] + MEM[7606];
assign MEM[35258] = MEM[7599] + MEM[7611];
assign MEM[35259] = MEM[7602] + MEM[7621];
assign MEM[35260] = MEM[7604] + MEM[7772];
assign MEM[35261] = MEM[7605] + MEM[8020];
assign MEM[35262] = MEM[7607] + MEM[7632];
assign MEM[35263] = MEM[7613] + MEM[7902];
assign MEM[35264] = MEM[7617] + MEM[7820];
assign MEM[35265] = MEM[7620] + MEM[7768];
assign MEM[35266] = MEM[7623] + MEM[8120];
assign MEM[35267] = MEM[7624] + MEM[7683];
assign MEM[35268] = MEM[7626] + MEM[7943];
assign MEM[35269] = MEM[7627] + MEM[7722];
assign MEM[35270] = MEM[7630] + MEM[7945];
assign MEM[35271] = MEM[7631] + MEM[7730];
assign MEM[35272] = MEM[7647] + MEM[7836];
assign MEM[35273] = MEM[7650] + MEM[7774];
assign MEM[35274] = MEM[7654] + MEM[7920];
assign MEM[35275] = MEM[7658] + MEM[7721];
assign MEM[35276] = MEM[7659] + MEM[7746];
assign MEM[35277] = MEM[7669] + MEM[7798];
assign MEM[35278] = MEM[7670] + MEM[7971];
assign MEM[35279] = MEM[7671] + MEM[7804];
assign MEM[35280] = MEM[7673] + MEM[7879];
assign MEM[35281] = MEM[7677] + MEM[7684];
assign MEM[35282] = MEM[7681] + MEM[8060];
assign MEM[35283] = MEM[7688] + MEM[7803];
assign MEM[35284] = MEM[7689] + MEM[7950];
assign MEM[35285] = MEM[7691] + MEM[7918];
assign MEM[35286] = MEM[7698] + MEM[7719];
assign MEM[35287] = MEM[7700] + MEM[7727];
assign MEM[35288] = MEM[7701] + MEM[7809];
assign MEM[35289] = MEM[7704] + MEM[7709];
assign MEM[35290] = MEM[7710] + MEM[7828];
assign MEM[35291] = MEM[7717] + MEM[7756];
assign MEM[35292] = MEM[7731] + MEM[7904];
assign MEM[35293] = MEM[7735] + MEM[7780];
assign MEM[35294] = MEM[7736] + MEM[7743];
assign MEM[35295] = MEM[7745] + MEM[7790];
assign MEM[35296] = MEM[7749] + MEM[7866];
assign MEM[35297] = MEM[7759] + MEM[7917];
assign MEM[35298] = MEM[7765] + MEM[7961];
assign MEM[35299] = MEM[7771] + MEM[7931];
assign MEM[35300] = MEM[7773] + MEM[7948];
assign MEM[35301] = MEM[7781] + MEM[8043];
assign MEM[35302] = MEM[7782] + MEM[7843];
assign MEM[35303] = MEM[7783] + MEM[7792];
assign MEM[35304] = MEM[7784] + MEM[7805];
assign MEM[35305] = MEM[7785] + MEM[7824];
assign MEM[35306] = MEM[7787] + MEM[7812];
assign MEM[35307] = MEM[7788] + MEM[8186];
assign MEM[35308] = MEM[7789] + MEM[7869];
assign MEM[35309] = MEM[7791] + MEM[7897];
assign MEM[35310] = MEM[7810] + MEM[7862];
assign MEM[35311] = MEM[7811] + MEM[7827];
assign MEM[35312] = MEM[7817] + MEM[7932];
assign MEM[35313] = MEM[7818] + MEM[7942];
assign MEM[35314] = MEM[7819] + MEM[7884];
assign MEM[35315] = MEM[7825] + MEM[8163];
assign MEM[35316] = MEM[7826] + MEM[7870];
assign MEM[35317] = MEM[7835] + MEM[7874];
assign MEM[35318] = MEM[7838] + MEM[7923];
assign MEM[35319] = MEM[7842] + MEM[7964];
assign MEM[35320] = MEM[7844] + MEM[8010];
assign MEM[35321] = MEM[7846] + MEM[7858];
assign MEM[35322] = MEM[7851] + MEM[7852];
assign MEM[35323] = MEM[7854] + MEM[8015];
assign MEM[35324] = MEM[7860] + MEM[7873];
assign MEM[35325] = MEM[7868] + MEM[8096];
assign MEM[35326] = MEM[7875] + MEM[8008];
assign MEM[35327] = MEM[7887] + MEM[7913];
assign MEM[35328] = MEM[7889] + MEM[7940];
assign MEM[35329] = MEM[7891] + MEM[7925];
assign MEM[35330] = MEM[7892] + MEM[7939];
assign MEM[35331] = MEM[7898] + MEM[7965];
assign MEM[35332] = MEM[7900] + MEM[8078];
assign MEM[35333] = MEM[7901] + MEM[8052];
assign MEM[35334] = MEM[7903] + MEM[8085];
assign MEM[35335] = MEM[7912] + MEM[7974];
assign MEM[35336] = MEM[7919] + MEM[7957];
assign MEM[35337] = MEM[7926] + MEM[8212];
assign MEM[35338] = MEM[7928] + MEM[8013];
assign MEM[35339] = MEM[7937] + MEM[8123];
assign MEM[35340] = MEM[7941] + MEM[8081];
assign MEM[35341] = MEM[7947] + MEM[8162];
assign MEM[35342] = MEM[7952] + MEM[8297];
assign MEM[35343] = MEM[7956] + MEM[8231];
assign MEM[35344] = MEM[7958] + MEM[7989];
assign MEM[35345] = MEM[7960] + MEM[7982];
assign MEM[35346] = MEM[7962] + MEM[7995];
assign MEM[35347] = MEM[7967] + MEM[8176];
assign MEM[35348] = MEM[7968] + MEM[8319];
assign MEM[35349] = MEM[7969] + MEM[8025];
assign MEM[35350] = MEM[7976] + MEM[8199];
assign MEM[35351] = MEM[7981] + MEM[8050];
assign MEM[35352] = MEM[7983] + MEM[8011];
assign MEM[35353] = MEM[7984] + MEM[8098];
assign MEM[35354] = MEM[7988] + MEM[8068];
assign MEM[35355] = MEM[7992] + MEM[8239];
assign MEM[35356] = MEM[7997] + MEM[8108];
assign MEM[35357] = MEM[8003] + MEM[8082];
assign MEM[35358] = MEM[8004] + MEM[8076];
assign MEM[35359] = MEM[8012] + MEM[8214];
assign MEM[35360] = MEM[8017] + MEM[8061];
assign MEM[35361] = MEM[8021] + MEM[8117];
assign MEM[35362] = MEM[8024] + MEM[8220];
assign MEM[35363] = MEM[8026] + MEM[8056];
assign MEM[35364] = MEM[8027] + MEM[8111];
assign MEM[35365] = MEM[8029] + MEM[8304];
assign MEM[35366] = MEM[8030] + MEM[8149];
assign MEM[35367] = MEM[8031] + MEM[8191];
assign MEM[35368] = MEM[8033] + MEM[8409];
assign MEM[35369] = MEM[8034] + MEM[8058];
assign MEM[35370] = MEM[8035] + MEM[8141];
assign MEM[35371] = MEM[8037] + MEM[8065];
assign MEM[35372] = MEM[8038] + MEM[8062];
assign MEM[35373] = MEM[8044] + MEM[8452];
assign MEM[35374] = MEM[8045] + MEM[8222];
assign MEM[35375] = MEM[8049] + MEM[8088];
assign MEM[35376] = MEM[8054] + MEM[8160];
assign MEM[35377] = MEM[8064] + MEM[8127];
assign MEM[35378] = MEM[8066] + MEM[8211];
assign MEM[35379] = MEM[8074] + MEM[8221];
assign MEM[35380] = MEM[8077] + MEM[8269];
assign MEM[35381] = MEM[8083] + MEM[8366];
assign MEM[35382] = MEM[8086] + MEM[8185];
assign MEM[35383] = MEM[8087] + MEM[8159];
assign MEM[35384] = MEM[8104] + MEM[8436];
assign MEM[35385] = MEM[8105] + MEM[8339];
assign MEM[35386] = MEM[8106] + MEM[8401];
assign MEM[35387] = MEM[8112] + MEM[8140];
assign MEM[35388] = MEM[8115] + MEM[8175];
assign MEM[35389] = MEM[8118] + MEM[8329];
assign MEM[35390] = MEM[8121] + MEM[8286];
assign MEM[35391] = MEM[8124] + MEM[8201];
assign MEM[35392] = MEM[8126] + MEM[8515];
assign MEM[35393] = MEM[8128] + MEM[8203];
assign MEM[35394] = MEM[8131] + MEM[8241];
assign MEM[35395] = MEM[8137] + MEM[8225];
assign MEM[35396] = MEM[8138] + MEM[8281];
assign MEM[35397] = MEM[8139] + MEM[8307];
assign MEM[35398] = MEM[8146] + MEM[8182];
assign MEM[35399] = MEM[8165] + MEM[8205];
assign MEM[35400] = MEM[8166] + MEM[8402];
assign MEM[35401] = MEM[8167] + MEM[8262];
assign MEM[35402] = MEM[8172] + MEM[8450];
assign MEM[35403] = MEM[8188] + MEM[8479];
assign MEM[35404] = MEM[8190] + MEM[8532];
assign MEM[35405] = MEM[8193] + MEM[8234];
assign MEM[35406] = MEM[8208] + MEM[8291];
assign MEM[35407] = MEM[8209] + MEM[8303];
assign MEM[35408] = MEM[8217] + MEM[8253];
assign MEM[35409] = MEM[8224] + MEM[8277];
assign MEM[35410] = MEM[8227] + MEM[8487];
assign MEM[35411] = MEM[8228] + MEM[8309];
assign MEM[35412] = MEM[8232] + MEM[8383];
assign MEM[35413] = MEM[8236] + MEM[8287];
assign MEM[35414] = MEM[8242] + MEM[8482];
assign MEM[35415] = MEM[8244] + MEM[8246];
assign MEM[35416] = MEM[8245] + MEM[8323];
assign MEM[35417] = MEM[8250] + MEM[8256];
assign MEM[35418] = MEM[8251] + MEM[8596];
assign MEM[35419] = MEM[8254] + MEM[8335];
assign MEM[35420] = MEM[8264] + MEM[8289];
assign MEM[35421] = MEM[8268] + MEM[8348];
assign MEM[35422] = MEM[8272] + MEM[8395];
assign MEM[35423] = MEM[8275] + MEM[8315];
assign MEM[35424] = MEM[8284] + MEM[8413];
assign MEM[35425] = MEM[8290] + MEM[8311];
assign MEM[35426] = MEM[8292] + MEM[8338];
assign MEM[35427] = MEM[8293] + MEM[8465];
assign MEM[35428] = MEM[8296] + MEM[8429];
assign MEM[35429] = MEM[8299] + MEM[8354];
assign MEM[35430] = MEM[8301] + MEM[8367];
assign MEM[35431] = MEM[8305] + MEM[8306];
assign MEM[35432] = MEM[8308] + MEM[8314];
assign MEM[35433] = MEM[8312] + MEM[8403];
assign MEM[35434] = MEM[8313] + MEM[8410];
assign MEM[35435] = MEM[8317] + MEM[8387];
assign MEM[35436] = MEM[8327] + MEM[8390];
assign MEM[35437] = MEM[8332] + MEM[8388];
assign MEM[35438] = MEM[8333] + MEM[8588];
assign MEM[35439] = MEM[8336] + MEM[8346];
assign MEM[35440] = MEM[8344] + MEM[8407];
assign MEM[35441] = MEM[8349] + MEM[8470];
assign MEM[35442] = MEM[8352] + MEM[8358];
assign MEM[35443] = MEM[8353] + MEM[8363];
assign MEM[35444] = MEM[8357] + MEM[8555];
assign MEM[35445] = MEM[8362] + MEM[8706];
assign MEM[35446] = MEM[8364] + MEM[8463];
assign MEM[35447] = MEM[8370] + MEM[8663];
assign MEM[35448] = MEM[8372] + MEM[8394];
assign MEM[35449] = MEM[8384] + MEM[8484];
assign MEM[35450] = MEM[8386] + MEM[8711];
assign MEM[35451] = MEM[8391] + MEM[8530];
assign MEM[35452] = MEM[8393] + MEM[8538];
assign MEM[35453] = MEM[8398] + MEM[8444];
assign MEM[35454] = MEM[8404] + MEM[8458];
assign MEM[35455] = MEM[8406] + MEM[8512];
assign MEM[35456] = MEM[8408] + MEM[8528];
assign MEM[35457] = MEM[8411] + MEM[8559];
assign MEM[35458] = MEM[8419] + MEM[8478];
assign MEM[35459] = MEM[8420] + MEM[8525];
assign MEM[35460] = MEM[8424] + MEM[8472];
assign MEM[35461] = MEM[8432] + MEM[8491];
assign MEM[35462] = MEM[8437] + MEM[8799];
assign MEM[35463] = MEM[8441] + MEM[8456];
assign MEM[35464] = MEM[8447] + MEM[8475];
assign MEM[35465] = MEM[8451] + MEM[8468];
assign MEM[35466] = MEM[8459] + MEM[8700];
assign MEM[35467] = MEM[8460] + MEM[8518];
assign MEM[35468] = MEM[8462] + MEM[8519];
assign MEM[35469] = MEM[8464] + MEM[8485];
assign MEM[35470] = MEM[8474] + MEM[8767];
assign MEM[35471] = MEM[8480] + MEM[8537];
assign MEM[35472] = MEM[8481] + MEM[8583];
assign MEM[35473] = MEM[8488] + MEM[8506];
assign MEM[35474] = MEM[8494] + MEM[8553];
assign MEM[35475] = MEM[8500] + MEM[8657];
assign MEM[35476] = MEM[8502] + MEM[8533];
assign MEM[35477] = MEM[8509] + MEM[8554];
assign MEM[35478] = MEM[8511] + MEM[8661];
assign MEM[35479] = MEM[8524] + MEM[8568];
assign MEM[35480] = MEM[8529] + MEM[8573];
assign MEM[35481] = MEM[8531] + MEM[8641];
assign MEM[35482] = MEM[8536] + MEM[8823];
assign MEM[35483] = MEM[8539] + MEM[8548];
assign MEM[35484] = MEM[8540] + MEM[8577];
assign MEM[35485] = MEM[8542] + MEM[9158];
assign MEM[35486] = MEM[8543] + MEM[8736];
assign MEM[35487] = MEM[8544] + MEM[8597];
assign MEM[35488] = MEM[8549] + MEM[8611];
assign MEM[35489] = MEM[8550] + MEM[8584];
assign MEM[35490] = MEM[8551] + MEM[8609];
assign MEM[35491] = MEM[8562] + MEM[8659];
assign MEM[35492] = MEM[8569] + MEM[8779];
assign MEM[35493] = MEM[8575] + MEM[8752];
assign MEM[35494] = MEM[8576] + MEM[8710];
assign MEM[35495] = MEM[8578] + MEM[8601];
assign MEM[35496] = MEM[8579] + MEM[8645];
assign MEM[35497] = MEM[8582] + MEM[8640];
assign MEM[35498] = MEM[8591] + MEM[8619];
assign MEM[35499] = MEM[8595] + MEM[8603];
assign MEM[35500] = MEM[8599] + MEM[8898];
assign MEM[35501] = MEM[8605] + MEM[8713];
assign MEM[35502] = MEM[8610] + MEM[8694];
assign MEM[35503] = MEM[8614] + MEM[8793];
assign MEM[35504] = MEM[8616] + MEM[8766];
assign MEM[35505] = MEM[8630] + MEM[8744];
assign MEM[35506] = MEM[8638] + MEM[8642];
assign MEM[35507] = MEM[8644] + MEM[8708];
assign MEM[35508] = MEM[8646] + MEM[8727];
assign MEM[35509] = MEM[8650] + MEM[8673];
assign MEM[35510] = MEM[8651] + MEM[8743];
assign MEM[35511] = MEM[8653] + MEM[8707];
assign MEM[35512] = MEM[8655] + MEM[8689];
assign MEM[35513] = MEM[8662] + MEM[8664];
assign MEM[35514] = MEM[8665] + MEM[8829];
assign MEM[35515] = MEM[8672] + MEM[8717];
assign MEM[35516] = MEM[8675] + MEM[8686];
assign MEM[35517] = MEM[8681] + MEM[9078];
assign MEM[35518] = MEM[8684] + MEM[8941];
assign MEM[35519] = MEM[8685] + MEM[8789];
assign MEM[35520] = MEM[8687] + MEM[8810];
assign MEM[35521] = MEM[8688] + MEM[9531];
assign MEM[35522] = MEM[8690] + MEM[9109];
assign MEM[35523] = MEM[8695] + MEM[8803];
assign MEM[35524] = MEM[8698] + MEM[8903];
assign MEM[35525] = MEM[8714] + MEM[8725];
assign MEM[35526] = MEM[8715] + MEM[8919];
assign MEM[35527] = MEM[8716] + MEM[8853];
assign MEM[35528] = MEM[8718] + MEM[8999];
assign MEM[35529] = MEM[8719] + MEM[8780];
assign MEM[35530] = MEM[8720] + MEM[8831];
assign MEM[35531] = MEM[8723] + MEM[8913];
assign MEM[35532] = MEM[8724] + MEM[8819];
assign MEM[35533] = MEM[8729] + MEM[8730];
assign MEM[35534] = MEM[8741] + MEM[8970];
assign MEM[35535] = MEM[8745] + MEM[9155];
assign MEM[35536] = MEM[8749] + MEM[8885];
assign MEM[35537] = MEM[8754] + MEM[8760];
assign MEM[35538] = MEM[8755] + MEM[9000];
assign MEM[35539] = MEM[8758] + MEM[8817];
assign MEM[35540] = MEM[8761] + MEM[8850];
assign MEM[35541] = MEM[8765] + MEM[8786];
assign MEM[35542] = MEM[8771] + MEM[8976];
assign MEM[35543] = MEM[8772] + MEM[8917];
assign MEM[35544] = MEM[8775] + MEM[9042];
assign MEM[35545] = MEM[8783] + MEM[8838];
assign MEM[35546] = MEM[8785] + MEM[8878];
assign MEM[35547] = MEM[8787] + MEM[8902];
assign MEM[35548] = MEM[8790] + MEM[8796];
assign MEM[35549] = MEM[8791] + MEM[8899];
assign MEM[35550] = MEM[8800] + MEM[8905];
assign MEM[35551] = MEM[8806] + MEM[8818];
assign MEM[35552] = MEM[8812] + MEM[8824];
assign MEM[35553] = MEM[8821] + MEM[8828];
assign MEM[35554] = MEM[8822] + MEM[8944];
assign MEM[35555] = MEM[8834] + MEM[9193];
assign MEM[35556] = MEM[8843] + MEM[8873];
assign MEM[35557] = MEM[8845] + MEM[9001];
assign MEM[35558] = MEM[8846] + MEM[8865];
assign MEM[35559] = MEM[8847] + MEM[9044];
assign MEM[35560] = MEM[8849] + MEM[9062];
assign MEM[35561] = MEM[8857] + MEM[8900];
assign MEM[35562] = MEM[8859] + MEM[8872];
assign MEM[35563] = MEM[8862] + MEM[9151];
assign MEM[35564] = MEM[8866] + MEM[9005];
assign MEM[35565] = MEM[8870] + MEM[8881];
assign MEM[35566] = MEM[8877] + MEM[8932];
assign MEM[35567] = MEM[8879] + MEM[9056];
assign MEM[35568] = MEM[8880] + MEM[9053];
assign MEM[35569] = MEM[8883] + MEM[8933];
assign MEM[35570] = MEM[8884] + MEM[9150];
assign MEM[35571] = MEM[8886] + MEM[9002];
assign MEM[35572] = MEM[8897] + MEM[8948];
assign MEM[35573] = MEM[8904] + MEM[8991];
assign MEM[35574] = MEM[8908] + MEM[9286];
assign MEM[35575] = MEM[8909] + MEM[9055];
assign MEM[35576] = MEM[8911] + MEM[9077];
assign MEM[35577] = MEM[8914] + MEM[9110];
assign MEM[35578] = MEM[8915] + MEM[9073];
assign MEM[35579] = MEM[8916] + MEM[8962];
assign MEM[35580] = MEM[8918] + MEM[9054];
assign MEM[35581] = MEM[8920] + MEM[9017];
assign MEM[35582] = MEM[8922] + MEM[9197];
assign MEM[35583] = MEM[8923] + MEM[9085];
assign MEM[35584] = MEM[8924] + MEM[9016];
assign MEM[35585] = MEM[8930] + MEM[8990];
assign MEM[35586] = MEM[8935] + MEM[8942];
assign MEM[35587] = MEM[8936] + MEM[9067];
assign MEM[35588] = MEM[8940] + MEM[8985];
assign MEM[35589] = MEM[8943] + MEM[8981];
assign MEM[35590] = MEM[8947] + MEM[9178];
assign MEM[35591] = MEM[8952] + MEM[9012];
assign MEM[35592] = MEM[8953] + MEM[9381];
assign MEM[35593] = MEM[8954] + MEM[8978];
assign MEM[35594] = MEM[8956] + MEM[9172];
assign MEM[35595] = MEM[8958] + MEM[9009];
assign MEM[35596] = MEM[8963] + MEM[9014];
assign MEM[35597] = MEM[8968] + MEM[9097];
assign MEM[35598] = MEM[8987] + MEM[9160];
assign MEM[35599] = MEM[8988] + MEM[9136];
assign MEM[35600] = MEM[8989] + MEM[9021];
assign MEM[35601] = MEM[8993] + MEM[9029];
assign MEM[35602] = MEM[8995] + MEM[9130];
assign MEM[35603] = MEM[9007] + MEM[9025];
assign MEM[35604] = MEM[9024] + MEM[9452];
assign MEM[35605] = MEM[9026] + MEM[9098];
assign MEM[35606] = MEM[9030] + MEM[9138];
assign MEM[35607] = MEM[9031] + MEM[9247];
assign MEM[35608] = MEM[9032] + MEM[9147];
assign MEM[35609] = MEM[9033] + MEM[9149];
assign MEM[35610] = MEM[9036] + MEM[9112];
assign MEM[35611] = MEM[9043] + MEM[9552];
assign MEM[35612] = MEM[9045] + MEM[9050];
assign MEM[35613] = MEM[9046] + MEM[9133];
assign MEM[35614] = MEM[9052] + MEM[9216];
assign MEM[35615] = MEM[9058] + MEM[9093];
assign MEM[35616] = MEM[9059] + MEM[9305];
assign MEM[35617] = MEM[9061] + MEM[9065];
assign MEM[35618] = MEM[9063] + MEM[9096];
assign MEM[35619] = MEM[9071] + MEM[9182];
assign MEM[35620] = MEM[9075] + MEM[9108];
assign MEM[35621] = MEM[9076] + MEM[9102];
assign MEM[35622] = MEM[9081] + MEM[9094];
assign MEM[35623] = MEM[9082] + MEM[9118];
assign MEM[35624] = MEM[9090] + MEM[9238];
assign MEM[35625] = MEM[9095] + MEM[9497];
assign MEM[35626] = MEM[9099] + MEM[9123];
assign MEM[35627] = MEM[9100] + MEM[9116];
assign MEM[35628] = MEM[9101] + MEM[9154];
assign MEM[35629] = MEM[9104] + MEM[9156];
assign MEM[35630] = MEM[9106] + MEM[9744];
assign MEM[35631] = MEM[9107] + MEM[9127];
assign MEM[35632] = MEM[9111] + MEM[9276];
assign MEM[35633] = MEM[9113] + MEM[9386];
assign MEM[35634] = MEM[9117] + MEM[9234];
assign MEM[35635] = MEM[9119] + MEM[9240];
assign MEM[35636] = MEM[9122] + MEM[9180];
assign MEM[35637] = MEM[9126] + MEM[9222];
assign MEM[35638] = MEM[9129] + MEM[9140];
assign MEM[35639] = MEM[9131] + MEM[9202];
assign MEM[35640] = MEM[9134] + MEM[9186];
assign MEM[35641] = MEM[9141] + MEM[9322];
assign MEM[35642] = MEM[9143] + MEM[9215];
assign MEM[35643] = MEM[9146] + MEM[9559];
assign MEM[35644] = MEM[9152] + MEM[9170];
assign MEM[35645] = MEM[9153] + MEM[9337];
assign MEM[35646] = MEM[9157] + MEM[9236];
assign MEM[35647] = MEM[9159] + MEM[9251];
assign MEM[35648] = MEM[9161] + MEM[9342];
assign MEM[35649] = MEM[9167] + MEM[9235];
assign MEM[35650] = MEM[9168] + MEM[9300];
assign MEM[35651] = MEM[9171] + MEM[9445];
assign MEM[35652] = MEM[9174] + MEM[9181];
assign MEM[35653] = MEM[9177] + MEM[9199];
assign MEM[35654] = MEM[9179] + MEM[9253];
assign MEM[35655] = MEM[9188] + MEM[9230];
assign MEM[35656] = MEM[9191] + MEM[9223];
assign MEM[35657] = MEM[9198] + MEM[9285];
assign MEM[35658] = MEM[9200] + MEM[9207];
assign MEM[35659] = MEM[9203] + MEM[9507];
assign MEM[35660] = MEM[9204] + MEM[9340];
assign MEM[35661] = MEM[9211] + MEM[9329];
assign MEM[35662] = MEM[9212] + MEM[9239];
assign MEM[35663] = MEM[9213] + MEM[9288];
assign MEM[35664] = MEM[9219] + MEM[9272];
assign MEM[35665] = MEM[9220] + MEM[9360];
assign MEM[35666] = MEM[9224] + MEM[9270];
assign MEM[35667] = MEM[9228] + MEM[9255];
assign MEM[35668] = MEM[9229] + MEM[9359];
assign MEM[35669] = MEM[9233] + MEM[9695];
assign MEM[35670] = MEM[9244] + MEM[9297];
assign MEM[35671] = MEM[9246] + MEM[9362];
assign MEM[35672] = MEM[9248] + MEM[9411];
assign MEM[35673] = MEM[9249] + MEM[9681];
assign MEM[35674] = MEM[9252] + MEM[9414];
assign MEM[35675] = MEM[9254] + MEM[9385];
assign MEM[35676] = MEM[9258] + MEM[9361];
assign MEM[35677] = MEM[9261] + MEM[9274];
assign MEM[35678] = MEM[9263] + MEM[9328];
assign MEM[35679] = MEM[9265] + MEM[9511];
assign MEM[35680] = MEM[9267] + MEM[9393];
assign MEM[35681] = MEM[9271] + MEM[9316];
assign MEM[35682] = MEM[9281] + MEM[9291];
assign MEM[35683] = MEM[9283] + MEM[9376];
assign MEM[35684] = MEM[9293] + MEM[9343];
assign MEM[35685] = MEM[9295] + MEM[9374];
assign MEM[35686] = MEM[9301] + MEM[9336];
assign MEM[35687] = MEM[9302] + MEM[9339];
assign MEM[35688] = MEM[9307] + MEM[9449];
assign MEM[35689] = MEM[9308] + MEM[9338];
assign MEM[35690] = MEM[9314] + MEM[9321];
assign MEM[35691] = MEM[9315] + MEM[9364];
assign MEM[35692] = MEM[9319] + MEM[9409];
assign MEM[35693] = MEM[9323] + MEM[9377];
assign MEM[35694] = MEM[9325] + MEM[9352];
assign MEM[35695] = MEM[9326] + MEM[9423];
assign MEM[35696] = MEM[9327] + MEM[9540];
assign MEM[35697] = MEM[9332] + MEM[9509];
assign MEM[35698] = MEM[9335] + MEM[9421];
assign MEM[35699] = MEM[9345] + MEM[9592];
assign MEM[35700] = MEM[9347] + MEM[9410];
assign MEM[35701] = MEM[9348] + MEM[9481];
assign MEM[35702] = MEM[9349] + MEM[9404];
assign MEM[35703] = MEM[9351] + MEM[9358];
assign MEM[35704] = MEM[9363] + MEM[9402];
assign MEM[35705] = MEM[9366] + MEM[9528];
assign MEM[35706] = MEM[9367] + MEM[9387];
assign MEM[35707] = MEM[9369] + MEM[9390];
assign MEM[35708] = MEM[9375] + MEM[9479];
assign MEM[35709] = MEM[9378] + MEM[9464];
assign MEM[35710] = MEM[9379] + MEM[9405];
assign MEM[35711] = MEM[9380] + MEM[9564];
assign MEM[35712] = MEM[9388] + MEM[9396];
assign MEM[35713] = MEM[9397] + MEM[9459];
assign MEM[35714] = MEM[9398] + MEM[9401];
assign MEM[35715] = MEM[9403] + MEM[9642];
assign MEM[35716] = MEM[9412] + MEM[9576];
assign MEM[35717] = MEM[9415] + MEM[9489];
assign MEM[35718] = MEM[9416] + MEM[9482];
assign MEM[35719] = MEM[9418] + MEM[9800];
assign MEM[35720] = MEM[9420] + MEM[9493];
assign MEM[35721] = MEM[9422] + MEM[9447];
assign MEM[35722] = MEM[9425] + MEM[9433];
assign MEM[35723] = MEM[9427] + MEM[9465];
assign MEM[35724] = MEM[9432] + MEM[9441];
assign MEM[35725] = MEM[9434] + MEM[9435];
assign MEM[35726] = MEM[9436] + MEM[9605];
assign MEM[35727] = MEM[9446] + MEM[9596];
assign MEM[35728] = MEM[9455] + MEM[9954];
assign MEM[35729] = MEM[9456] + MEM[9578];
assign MEM[35730] = MEM[9460] + MEM[9524];
assign MEM[35731] = MEM[9461] + MEM[9483];
assign MEM[35732] = MEM[9467] + MEM[9634];
assign MEM[35733] = MEM[9471] + MEM[9508];
assign MEM[35734] = MEM[9472] + MEM[9568];
assign MEM[35735] = MEM[9474] + MEM[9514];
assign MEM[35736] = MEM[9475] + MEM[9766];
assign MEM[35737] = MEM[9477] + MEM[9590];
assign MEM[35738] = MEM[9480] + MEM[9573];
assign MEM[35739] = MEM[9484] + MEM[9871];
assign MEM[35740] = MEM[9485] + MEM[9490];
assign MEM[35741] = MEM[9487] + MEM[9594];
assign MEM[35742] = MEM[9491] + MEM[9601];
assign MEM[35743] = MEM[9500] + MEM[9521];
assign MEM[35744] = MEM[9501] + MEM[9611];
assign MEM[35745] = MEM[9504] + MEM[9547];
assign MEM[35746] = MEM[9513] + MEM[9515];
assign MEM[35747] = MEM[9517] + MEM[9593];
assign MEM[35748] = MEM[9519] + MEM[9725];
assign MEM[35749] = MEM[9526] + MEM[9775];
assign MEM[35750] = MEM[9534] + MEM[9660];
assign MEM[35751] = MEM[9535] + MEM[9731];
assign MEM[35752] = MEM[9536] + MEM[9662];
assign MEM[35753] = MEM[9537] + MEM[9678];
assign MEM[35754] = MEM[9542] + MEM[9556];
assign MEM[35755] = MEM[9543] + MEM[9942];
assign MEM[35756] = MEM[9545] + MEM[9587];
assign MEM[35757] = MEM[9546] + MEM[9558];
assign MEM[35758] = MEM[9548] + MEM[9845];
assign MEM[35759] = MEM[9553] + MEM[9733];
assign MEM[35760] = MEM[9565] + MEM[9600];
assign MEM[35761] = MEM[9566] + MEM[9629];
assign MEM[35762] = MEM[9569] + MEM[9571];
assign MEM[35763] = MEM[9572] + MEM[9604];
assign MEM[35764] = MEM[9574] + MEM[9575];
assign MEM[35765] = MEM[9579] + MEM[9854];
assign MEM[35766] = MEM[9580] + MEM[9616];
assign MEM[35767] = MEM[9581] + MEM[9595];
assign MEM[35768] = MEM[9583] + MEM[9589];
assign MEM[35769] = MEM[9585] + MEM[9682];
assign MEM[35770] = MEM[9597] + MEM[9620];
assign MEM[35771] = MEM[9599] + MEM[9609];
assign MEM[35772] = MEM[9603] + MEM[9653];
assign MEM[35773] = MEM[9607] + MEM[9618];
assign MEM[35774] = MEM[9608] + MEM[9687];
assign MEM[35775] = MEM[9613] + MEM[9669];
assign MEM[35776] = MEM[9619] + MEM[9721];
assign MEM[35777] = MEM[9621] + MEM[10324];
assign MEM[35778] = MEM[9622] + MEM[9903];
assign MEM[35779] = MEM[9624] + MEM[9647];
assign MEM[35780] = MEM[9626] + MEM[9639];
assign MEM[35781] = MEM[9631] + MEM[9649];
assign MEM[35782] = MEM[9633] + MEM[9699];
assign MEM[35783] = MEM[9638] + MEM[9685];
assign MEM[35784] = MEM[9654] + MEM[9667];
assign MEM[35785] = MEM[9656] + MEM[9730];
assign MEM[35786] = MEM[9658] + MEM[9937];
assign MEM[35787] = MEM[9659] + MEM[9821];
assign MEM[35788] = MEM[9663] + MEM[9874];
assign MEM[35789] = MEM[9665] + MEM[9819];
assign MEM[35790] = MEM[9666] + MEM[9668];
assign MEM[35791] = MEM[9676] + MEM[9704];
assign MEM[35792] = MEM[9677] + MEM[9746];
assign MEM[35793] = MEM[9680] + MEM[9703];
assign MEM[35794] = MEM[9684] + MEM[9761];
assign MEM[35795] = MEM[9688] + MEM[9808];
assign MEM[35796] = MEM[9689] + MEM[9693];
assign MEM[35797] = MEM[9692] + MEM[9790];
assign MEM[35798] = MEM[9696] + MEM[9715];
assign MEM[35799] = MEM[9697] + MEM[10481];
assign MEM[35800] = MEM[9701] + MEM[9751];
assign MEM[35801] = MEM[9702] + MEM[9711];
assign MEM[35802] = MEM[9707] + MEM[9984];
assign MEM[35803] = MEM[9708] + MEM[10112];
assign MEM[35804] = MEM[9710] + MEM[9774];
assign MEM[35805] = MEM[9712] + MEM[9836];
assign MEM[35806] = MEM[9714] + MEM[10144];
assign MEM[35807] = MEM[9716] + MEM[10270];
assign MEM[35808] = MEM[9718] + MEM[9811];
assign MEM[35809] = MEM[9723] + MEM[9863];
assign MEM[35810] = MEM[9732] + MEM[9882];
assign MEM[35811] = MEM[9734] + MEM[10029];
assign MEM[35812] = MEM[9735] + MEM[9743];
assign MEM[35813] = MEM[9737] + MEM[9762];
assign MEM[35814] = MEM[9739] + MEM[9827];
assign MEM[35815] = MEM[9745] + MEM[9802];
assign MEM[35816] = MEM[9747] + MEM[9772];
assign MEM[35817] = MEM[9749] + MEM[9785];
assign MEM[35818] = MEM[9752] + MEM[9756];
assign MEM[35819] = MEM[9759] + MEM[9834];
assign MEM[35820] = MEM[9760] + MEM[10347];
assign MEM[35821] = MEM[9764] + MEM[9904];
assign MEM[35822] = MEM[9768] + MEM[10011];
assign MEM[35823] = MEM[9770] + MEM[9870];
assign MEM[35824] = MEM[9776] + MEM[9804];
assign MEM[35825] = MEM[9778] + MEM[9983];
assign MEM[35826] = MEM[9779] + MEM[9886];
assign MEM[35827] = MEM[9786] + MEM[9843];
assign MEM[35828] = MEM[9787] + MEM[9867];
assign MEM[35829] = MEM[9789] + MEM[9920];
assign MEM[35830] = MEM[9792] + MEM[9793];
assign MEM[35831] = MEM[9795] + MEM[9977];
assign MEM[35832] = MEM[9797] + MEM[9853];
assign MEM[35833] = MEM[9806] + MEM[9831];
assign MEM[35834] = MEM[9807] + MEM[9994];
assign MEM[35835] = MEM[9809] + MEM[9847];
assign MEM[35836] = MEM[9810] + MEM[9952];
assign MEM[35837] = MEM[9815] + MEM[9859];
assign MEM[35838] = MEM[9818] + MEM[9926];
assign MEM[35839] = MEM[9828] + MEM[9855];
assign MEM[35840] = MEM[9829] + MEM[10303];
assign MEM[35841] = MEM[9832] + MEM[9951];
assign MEM[35842] = MEM[9833] + MEM[9868];
assign MEM[35843] = MEM[9837] + MEM[9950];
assign MEM[35844] = MEM[9838] + MEM[9940];
assign MEM[35845] = MEM[9842] + MEM[9915];
assign MEM[35846] = MEM[9844] + MEM[9948];
assign MEM[35847] = MEM[9846] + MEM[9932];
assign MEM[35848] = MEM[9849] + MEM[10058];
assign MEM[35849] = MEM[9850] + MEM[9999];
assign MEM[35850] = MEM[9852] + MEM[10026];
assign MEM[35851] = MEM[9858] + MEM[9936];
assign MEM[35852] = MEM[9865] + MEM[9928];
assign MEM[35853] = MEM[9873] + MEM[10152];
assign MEM[35854] = MEM[9876] + MEM[9911];
assign MEM[35855] = MEM[9878] + MEM[9916];
assign MEM[35856] = MEM[9880] + MEM[9914];
assign MEM[35857] = MEM[9883] + MEM[9890];
assign MEM[35858] = MEM[9892] + MEM[9995];
assign MEM[35859] = MEM[9895] + MEM[9996];
assign MEM[35860] = MEM[9905] + MEM[10010];
assign MEM[35861] = MEM[9906] + MEM[10285];
assign MEM[35862] = MEM[9909] + MEM[9927];
assign MEM[35863] = MEM[9910] + MEM[9912];
assign MEM[35864] = MEM[9913] + MEM[9933];
assign MEM[35865] = MEM[9917] + MEM[10163];
assign MEM[35866] = MEM[9919] + MEM[9960];
assign MEM[35867] = MEM[9922] + MEM[9931];
assign MEM[35868] = MEM[9929] + MEM[9968];
assign MEM[35869] = MEM[9934] + MEM[10214];
assign MEM[35870] = MEM[9935] + MEM[10051];
assign MEM[35871] = MEM[9938] + MEM[10043];
assign MEM[35872] = MEM[9939] + MEM[10033];
assign MEM[35873] = MEM[9941] + MEM[9961];
assign MEM[35874] = MEM[9949] + MEM[9989];
assign MEM[35875] = MEM[9955] + MEM[10042];
assign MEM[35876] = MEM[9956] + MEM[10065];
assign MEM[35877] = MEM[9958] + MEM[10053];
assign MEM[35878] = MEM[9966] + MEM[10119];
assign MEM[35879] = MEM[9972] + MEM[10121];
assign MEM[35880] = MEM[9973] + MEM[10003];
assign MEM[35881] = MEM[9975] + MEM[10031];
assign MEM[35882] = MEM[9978] + MEM[10049];
assign MEM[35883] = MEM[9986] + MEM[10077];
assign MEM[35884] = MEM[9990] + MEM[10113];
assign MEM[35885] = MEM[9991] + MEM[10179];
assign MEM[35886] = MEM[9992] + MEM[10025];
assign MEM[35887] = MEM[10005] + MEM[10022];
assign MEM[35888] = MEM[10007] + MEM[10019];
assign MEM[35889] = MEM[10008] + MEM[10068];
assign MEM[35890] = MEM[10009] + MEM[10229];
assign MEM[35891] = MEM[10012] + MEM[10452];
assign MEM[35892] = MEM[10013] + MEM[10255];
assign MEM[35893] = MEM[10015] + MEM[10032];
assign MEM[35894] = MEM[10016] + MEM[10020];
assign MEM[35895] = MEM[10018] + MEM[10050];
assign MEM[35896] = MEM[10027] + MEM[10189];
assign MEM[35897] = MEM[10039] + MEM[10066];
assign MEM[35898] = MEM[10040] + MEM[10160];
assign MEM[35899] = MEM[10041] + MEM[10317];
assign MEM[35900] = MEM[10046] + MEM[10370];
assign MEM[35901] = MEM[10048] + MEM[10353];
assign MEM[35902] = MEM[10054] + MEM[10106];
assign MEM[35903] = MEM[10057] + MEM[11383];
assign MEM[35904] = MEM[10060] + MEM[10171];
assign MEM[35905] = MEM[10061] + MEM[10072];
assign MEM[35906] = MEM[10071] + MEM[10169];
assign MEM[35907] = MEM[10074] + MEM[10086];
assign MEM[35908] = MEM[10081] + MEM[10126];
assign MEM[35909] = MEM[10087] + MEM[10276];
assign MEM[35910] = MEM[10088] + MEM[10166];
assign MEM[35911] = MEM[10091] + MEM[10129];
assign MEM[35912] = MEM[10092] + MEM[10192];
assign MEM[35913] = MEM[10105] + MEM[10200];
assign MEM[35914] = MEM[10111] + MEM[10142];
assign MEM[35915] = MEM[10114] + MEM[10157];
assign MEM[35916] = MEM[10115] + MEM[10258];
assign MEM[35917] = MEM[10118] + MEM[10161];
assign MEM[35918] = MEM[10127] + MEM[10268];
assign MEM[35919] = MEM[10131] + MEM[10320];
assign MEM[35920] = MEM[10135] + MEM[10244];
assign MEM[35921] = MEM[10137] + MEM[10150];
assign MEM[35922] = MEM[10138] + MEM[10170];
assign MEM[35923] = MEM[10145] + MEM[10260];
assign MEM[35924] = MEM[10146] + MEM[10318];
assign MEM[35925] = MEM[10149] + MEM[10273];
assign MEM[35926] = MEM[10154] + MEM[10158];
assign MEM[35927] = MEM[10155] + MEM[10223];
assign MEM[35928] = MEM[10162] + MEM[10194];
assign MEM[35929] = MEM[10165] + MEM[10291];
assign MEM[35930] = MEM[10167] + MEM[10186];
assign MEM[35931] = MEM[10168] + MEM[10206];
assign MEM[35932] = MEM[10180] + MEM[10522];
assign MEM[35933] = MEM[10184] + MEM[10434];
assign MEM[35934] = MEM[10188] + MEM[10362];
assign MEM[35935] = MEM[10196] + MEM[10226];
assign MEM[35936] = MEM[10199] + MEM[10212];
assign MEM[35937] = MEM[10202] + MEM[10267];
assign MEM[35938] = MEM[10204] + MEM[10333];
assign MEM[35939] = MEM[10207] + MEM[10314];
assign MEM[35940] = MEM[10209] + MEM[10221];
assign MEM[35941] = MEM[10210] + MEM[10589];
assign MEM[35942] = MEM[10211] + MEM[10520];
assign MEM[35943] = MEM[10215] + MEM[10339];
assign MEM[35944] = MEM[10222] + MEM[10366];
assign MEM[35945] = MEM[10230] + MEM[10483];
assign MEM[35946] = MEM[10237] + MEM[10490];
assign MEM[35947] = MEM[10239] + MEM[10287];
assign MEM[35948] = MEM[10243] + MEM[10252];
assign MEM[35949] = MEM[10245] + MEM[10567];
assign MEM[35950] = MEM[10259] + MEM[10281];
assign MEM[35951] = MEM[10264] + MEM[10295];
assign MEM[35952] = MEM[10274] + MEM[10348];
assign MEM[35953] = MEM[10275] + MEM[10449];
assign MEM[35954] = MEM[10282] + MEM[10354];
assign MEM[35955] = MEM[10284] + MEM[10462];
assign MEM[35956] = MEM[10290] + MEM[10473];
assign MEM[35957] = MEM[10294] + MEM[10479];
assign MEM[35958] = MEM[10296] + MEM[10430];
assign MEM[35959] = MEM[10297] + MEM[10443];
assign MEM[35960] = MEM[10299] + MEM[10529];
assign MEM[35961] = MEM[10300] + MEM[10380];
assign MEM[35962] = MEM[10306] + MEM[10402];
assign MEM[35963] = MEM[10307] + MEM[10786];
assign MEM[35964] = MEM[10315] + MEM[10432];
assign MEM[35965] = MEM[10323] + MEM[10525];
assign MEM[35966] = MEM[10332] + MEM[10394];
assign MEM[35967] = MEM[10336] + MEM[10337];
assign MEM[35968] = MEM[10342] + MEM[10439];
assign MEM[35969] = MEM[10345] + MEM[10476];
assign MEM[35970] = MEM[10346] + MEM[10519];
assign MEM[35971] = MEM[10350] + MEM[10368];
assign MEM[35972] = MEM[10351] + MEM[10826];
assign MEM[35973] = MEM[10352] + MEM[10399];
assign MEM[35974] = MEM[10359] + MEM[10396];
assign MEM[35975] = MEM[10360] + MEM[10466];
assign MEM[35976] = MEM[10367] + MEM[10556];
assign MEM[35977] = MEM[10371] + MEM[10463];
assign MEM[35978] = MEM[10372] + MEM[10545];
assign MEM[35979] = MEM[10375] + MEM[10702];
assign MEM[35980] = MEM[10377] + MEM[10532];
assign MEM[35981] = MEM[10381] + MEM[10388];
assign MEM[35982] = MEM[10386] + MEM[10470];
assign MEM[35983] = MEM[10389] + MEM[10405];
assign MEM[35984] = MEM[10398] + MEM[10477];
assign MEM[35985] = MEM[10400] + MEM[10537];
assign MEM[35986] = MEM[10401] + MEM[10631];
assign MEM[35987] = MEM[10406] + MEM[10726];
assign MEM[35988] = MEM[10409] + MEM[10559];
assign MEM[35989] = MEM[10410] + MEM[10448];
assign MEM[35990] = MEM[10417] + MEM[10760];
assign MEM[35991] = MEM[10418] + MEM[10586];
assign MEM[35992] = MEM[10431] + MEM[10446];
assign MEM[35993] = MEM[10433] + MEM[10534];
assign MEM[35994] = MEM[10451] + MEM[10461];
assign MEM[35995] = MEM[10464] + MEM[10632];
assign MEM[35996] = MEM[10467] + MEM[10510];
assign MEM[35997] = MEM[10468] + MEM[11246];
assign MEM[35998] = MEM[10478] + MEM[10856];
assign MEM[35999] = MEM[10482] + MEM[11072];
assign MEM[36000] = MEM[10492] + MEM[10541];
assign MEM[36001] = MEM[10506] + MEM[10721];
assign MEM[36002] = MEM[10507] + MEM[10944];
assign MEM[36003] = MEM[10508] + MEM[10705];
assign MEM[36004] = MEM[10516] + MEM[11182];
assign MEM[36005] = MEM[10518] + MEM[10718];
assign MEM[36006] = MEM[10523] + MEM[11301];
assign MEM[36007] = MEM[10531] + MEM[10637];
assign MEM[36008] = MEM[10536] + MEM[10692];
assign MEM[36009] = MEM[10549] + MEM[10554];
assign MEM[36010] = MEM[10557] + MEM[11034];
assign MEM[36011] = MEM[10558] + MEM[10840];
assign MEM[36012] = MEM[10560] + MEM[10751];
assign MEM[36013] = MEM[10573] + MEM[11008];
assign MEM[36014] = MEM[10578] + MEM[10640];
assign MEM[36015] = MEM[10581] + MEM[11025];
assign MEM[36016] = MEM[10593] + MEM[10894];
assign MEM[36017] = MEM[10596] + MEM[10605];
assign MEM[36018] = MEM[10600] + MEM[10765];
assign MEM[36019] = MEM[10608] + MEM[10615];
assign MEM[36020] = MEM[10609] + MEM[10794];
assign MEM[36021] = MEM[10611] + MEM[11146];
assign MEM[36022] = MEM[10619] + MEM[11340];
assign MEM[36023] = MEM[10620] + MEM[11286];
assign MEM[36024] = MEM[10634] + MEM[10995];
assign MEM[36025] = MEM[10638] + MEM[10708];
assign MEM[36026] = MEM[10643] + MEM[11099];
assign MEM[36027] = MEM[10644] + MEM[11019];
assign MEM[36028] = MEM[10656] + MEM[11031];
assign MEM[36029] = MEM[10659] + MEM[10912];
assign MEM[36030] = MEM[10662] + MEM[10703];
assign MEM[36031] = MEM[10664] + MEM[10752];
assign MEM[36032] = MEM[10675] + MEM[10891];
assign MEM[36033] = MEM[10681] + MEM[11196];
assign MEM[36034] = MEM[10684] + MEM[11027];
assign MEM[36035] = MEM[10685] + MEM[10727];
assign MEM[36036] = MEM[10699] + MEM[10924];
assign MEM[36037] = MEM[10716] + MEM[10887];
assign MEM[36038] = MEM[10723] + MEM[10843];
assign MEM[36039] = MEM[10728] + MEM[10890];
assign MEM[36040] = MEM[10729] + MEM[11197];
assign MEM[36041] = MEM[10730] + MEM[11180];
assign MEM[36042] = MEM[10741] + MEM[11184];
assign MEM[36043] = MEM[10742] + MEM[10755];
assign MEM[36044] = MEM[10743] + MEM[10774];
assign MEM[36045] = MEM[10754] + MEM[10758];
assign MEM[36046] = MEM[10764] + MEM[10785];
assign MEM[36047] = MEM[10767] + MEM[11234];
assign MEM[36048] = MEM[10776] + MEM[10853];
assign MEM[36049] = MEM[10783] + MEM[10862];
assign MEM[36050] = MEM[10811] + MEM[11044];
assign MEM[36051] = MEM[10813] + MEM[11268];
assign MEM[36052] = MEM[10827] + MEM[10916];
assign MEM[36053] = MEM[10841] + MEM[10962];
assign MEM[36054] = MEM[10861] + MEM[11094];
assign MEM[36055] = MEM[10870] + MEM[10967];
assign MEM[36056] = MEM[10875] + MEM[11250];
assign MEM[36057] = MEM[10882] + MEM[10906];
assign MEM[36058] = MEM[10886] + MEM[10913];
assign MEM[36059] = MEM[10908] + MEM[11104];
assign MEM[36060] = MEM[10909] + MEM[11201];
assign MEM[36061] = MEM[10915] + MEM[11092];
assign MEM[36062] = MEM[10923] + MEM[11038];
assign MEM[36063] = MEM[10927] + MEM[11108];
assign MEM[36064] = MEM[10929] + MEM[10994];
assign MEM[36065] = MEM[10931] + MEM[11086];
assign MEM[36066] = MEM[10932] + MEM[11263];
assign MEM[36067] = MEM[10938] + MEM[10945];
assign MEM[36068] = MEM[10941] + MEM[11021];
assign MEM[36069] = MEM[10951] + MEM[11107];
assign MEM[36070] = MEM[10954] + MEM[11122];
assign MEM[36071] = MEM[10960] + MEM[11191];
assign MEM[36072] = MEM[10969] + MEM[11165];
assign MEM[36073] = MEM[10983] + MEM[11033];
assign MEM[36074] = MEM[11002] + MEM[11415];
assign MEM[36075] = MEM[11006] + MEM[11097];
assign MEM[36076] = MEM[11011] + MEM[11269];
assign MEM[36077] = MEM[11013] + MEM[11317];
assign MEM[36078] = MEM[11036] + MEM[11111];
assign MEM[36079] = MEM[11039] + MEM[11259];
assign MEM[36080] = MEM[11043] + MEM[11285];
assign MEM[36081] = MEM[11045] + MEM[11135];
assign MEM[36082] = MEM[11051] + MEM[11479];
assign MEM[36083] = MEM[11058] + MEM[11207];
assign MEM[36084] = MEM[11066] + MEM[11120];
assign MEM[36085] = MEM[11071] + MEM[11295];
assign MEM[36086] = MEM[11074] + MEM[11085];
assign MEM[36087] = MEM[11081] + MEM[11434];
assign MEM[36088] = MEM[11095] + MEM[11209];
assign MEM[36089] = MEM[11100] + MEM[11175];
assign MEM[36090] = MEM[11103] + MEM[11216];
assign MEM[36091] = MEM[11131] + MEM[11408];
assign MEM[36092] = MEM[11133] + MEM[11319];
assign MEM[36093] = MEM[11155] + MEM[11239];
assign MEM[36094] = MEM[11162] + MEM[11364];
assign MEM[36095] = MEM[11166] + MEM[11260];
assign MEM[36096] = MEM[11168] + MEM[11388];
assign MEM[36097] = MEM[11169] + MEM[11344];
assign MEM[36098] = MEM[11188] + MEM[11232];
assign MEM[36099] = MEM[11189] + MEM[11206];
assign MEM[36100] = MEM[11194] + MEM[11252];
assign MEM[36101] = MEM[11198] + MEM[11202];
assign MEM[36102] = MEM[11199] + MEM[11314];
assign MEM[36103] = MEM[11200] + MEM[11428];
assign MEM[36104] = MEM[11211] + MEM[11272];
assign MEM[36105] = MEM[11224] + MEM[11243];
assign MEM[36106] = MEM[11227] + MEM[11289];
assign MEM[36107] = MEM[11230] + MEM[11281];
assign MEM[36108] = MEM[11235] + MEM[11423];
assign MEM[36109] = MEM[11236] + MEM[11399];
assign MEM[36110] = MEM[11240] + MEM[11283];
assign MEM[36111] = MEM[11241] + MEM[11251];
assign MEM[36112] = MEM[11242] + MEM[11432];
assign MEM[36113] = MEM[11244] + MEM[11311];
assign MEM[36114] = MEM[11245] + MEM[11247];
assign MEM[36115] = MEM[11257] + MEM[11271];
assign MEM[36116] = MEM[11262] + MEM[11270];
assign MEM[36117] = MEM[11267] + MEM[11378];
assign MEM[36118] = MEM[11277] + MEM[11365];
assign MEM[36119] = MEM[11279] + MEM[11337];
assign MEM[36120] = MEM[11287] + MEM[11313];
assign MEM[36121] = MEM[11288] + MEM[11386];
assign MEM[36122] = MEM[11298] + MEM[11452];
assign MEM[36123] = MEM[11303] + MEM[11600];
assign MEM[36124] = MEM[11316] + MEM[11437];
assign MEM[36125] = MEM[11322] + MEM[11377];
assign MEM[36126] = MEM[11324] + MEM[11347];
assign MEM[36127] = MEM[11325] + MEM[11416];
assign MEM[36128] = MEM[11329] + MEM[11392];
assign MEM[36129] = MEM[11335] + MEM[11389];
assign MEM[36130] = MEM[11336] + MEM[11387];
assign MEM[36131] = MEM[11339] + MEM[11361];
assign MEM[36132] = MEM[11342] + MEM[11357];
assign MEM[36133] = MEM[11343] + MEM[11356];
assign MEM[36134] = MEM[11346] + MEM[11374];
assign MEM[36135] = MEM[11349] + MEM[11537];
assign MEM[36136] = MEM[11350] + MEM[11366];
assign MEM[36137] = MEM[11352] + MEM[11410];
assign MEM[36138] = MEM[11353] + MEM[11390];
assign MEM[36139] = MEM[11359] + MEM[11424];
assign MEM[36140] = MEM[11360] + MEM[11376];
assign MEM[36141] = MEM[11362] + MEM[11488];
assign MEM[36142] = MEM[11367] + MEM[11522];
assign MEM[36143] = MEM[11368] + MEM[11373];
assign MEM[36144] = MEM[11371] + MEM[11444];
assign MEM[36145] = MEM[11372] + MEM[11429];
assign MEM[36146] = MEM[11379] + MEM[11384];
assign MEM[36147] = MEM[11382] + MEM[11433];
assign MEM[36148] = MEM[11385] + MEM[11513];
assign MEM[36149] = MEM[11391] + MEM[11435];
assign MEM[36150] = MEM[11393] + MEM[11453];
assign MEM[36151] = MEM[11394] + MEM[11496];
assign MEM[36152] = MEM[11396] + MEM[11450];
assign MEM[36153] = MEM[11397] + MEM[11481];
assign MEM[36154] = MEM[11400] + MEM[11512];
assign MEM[36155] = MEM[11401] + MEM[11625];
assign MEM[36156] = MEM[11402] + MEM[11622];
assign MEM[36157] = MEM[11404] + MEM[11499];
assign MEM[36158] = MEM[11405] + MEM[11409];
assign MEM[36159] = MEM[11407] + MEM[11480];
assign MEM[36160] = MEM[11413] + MEM[11486];
assign MEM[36161] = MEM[11417] + MEM[11455];
assign MEM[36162] = MEM[11418] + MEM[11448];
assign MEM[36163] = MEM[11419] + MEM[11436];
assign MEM[36164] = MEM[11420] + MEM[11460];
assign MEM[36165] = MEM[11425] + MEM[11530];
assign MEM[36166] = MEM[11426] + MEM[11516];
assign MEM[36167] = MEM[11430] + MEM[11482];
assign MEM[36168] = MEM[11438] + MEM[11520];
assign MEM[36169] = MEM[11441] + MEM[11446];
assign MEM[36170] = MEM[11442] + MEM[11672];
assign MEM[36171] = MEM[11449] + MEM[11469];
assign MEM[36172] = MEM[11454] + MEM[11515];
assign MEM[36173] = MEM[11457] + MEM[11687];
assign MEM[36174] = MEM[11458] + MEM[11631];
assign MEM[36175] = MEM[11459] + MEM[11990];
assign MEM[36176] = MEM[11461] + MEM[12143];
assign MEM[36177] = MEM[11462] + MEM[11518];
assign MEM[36178] = MEM[11464] + MEM[11472];
assign MEM[36179] = MEM[11466] + MEM[11507];
assign MEM[36180] = MEM[11468] + MEM[11476];
assign MEM[36181] = MEM[11471] + MEM[11997];
assign MEM[36182] = MEM[11474] + MEM[11519];
assign MEM[36183] = MEM[11475] + MEM[11502];
assign MEM[36184] = MEM[11478] + MEM[11595];
assign MEM[36185] = MEM[11491] + MEM[11744];
assign MEM[36186] = MEM[11492] + MEM[11511];
assign MEM[36187] = MEM[11493] + MEM[11547];
assign MEM[36188] = MEM[11495] + MEM[11647];
assign MEM[36189] = MEM[11497] + MEM[11517];
assign MEM[36190] = MEM[11498] + MEM[11646];
assign MEM[36191] = MEM[11500] + MEM[11632];
assign MEM[36192] = MEM[11501] + MEM[11832];
assign MEM[36193] = MEM[11503] + MEM[11715];
assign MEM[36194] = MEM[11504] + MEM[11614];
assign MEM[36195] = MEM[11506] + MEM[11601];
assign MEM[36196] = MEM[11509] + MEM[11567];
assign MEM[36197] = MEM[11521] + MEM[11780];
assign MEM[36198] = MEM[11523] + MEM[11565];
assign MEM[36199] = MEM[11524] + MEM[11658];
assign MEM[36200] = MEM[11525] + MEM[11579];
assign MEM[36201] = MEM[11534] + MEM[11628];
assign MEM[36202] = MEM[11539] + MEM[11676];
assign MEM[36203] = MEM[11541] + MEM[11545];
assign MEM[36204] = MEM[11544] + MEM[11581];
assign MEM[36205] = MEM[11548] + MEM[11613];
assign MEM[36206] = MEM[11551] + MEM[11797];
assign MEM[36207] = MEM[11552] + MEM[11867];
assign MEM[36208] = MEM[11554] + MEM[11587];
assign MEM[36209] = MEM[11556] + MEM[11609];
assign MEM[36210] = MEM[11557] + MEM[11666];
assign MEM[36211] = MEM[11559] + MEM[11845];
assign MEM[36212] = MEM[11562] + MEM[11730];
assign MEM[36213] = MEM[11570] + MEM[11684];
assign MEM[36214] = MEM[11572] + MEM[11685];
assign MEM[36215] = MEM[11573] + MEM[11596];
assign MEM[36216] = MEM[11574] + MEM[11735];
assign MEM[36217] = MEM[11577] + MEM[11621];
assign MEM[36218] = MEM[11588] + MEM[11616];
assign MEM[36219] = MEM[11599] + MEM[11677];
assign MEM[36220] = MEM[11602] + MEM[11624];
assign MEM[36221] = MEM[11608] + MEM[11790];
assign MEM[36222] = MEM[11610] + MEM[11692];
assign MEM[36223] = MEM[11612] + MEM[11627];
assign MEM[36224] = MEM[11615] + MEM[11630];
assign MEM[36225] = MEM[11618] + MEM[11640];
assign MEM[36226] = MEM[11629] + MEM[11663];
assign MEM[36227] = MEM[11633] + MEM[11916];
assign MEM[36228] = MEM[11634] + MEM[11876];
assign MEM[36229] = MEM[11639] + MEM[11662];
assign MEM[36230] = MEM[11642] + MEM[11743];
assign MEM[36231] = MEM[11643] + MEM[11775];
assign MEM[36232] = MEM[11644] + MEM[12006];
assign MEM[36233] = MEM[11653] + MEM[11966];
assign MEM[36234] = MEM[11655] + MEM[11697];
assign MEM[36235] = MEM[11668] + MEM[11675];
assign MEM[36236] = MEM[11669] + MEM[11700];
assign MEM[36237] = MEM[11670] + MEM[11690];
assign MEM[36238] = MEM[11671] + MEM[11751];
assign MEM[36239] = MEM[11673] + MEM[11805];
assign MEM[36240] = MEM[11679] + MEM[11925];
assign MEM[36241] = MEM[11686] + MEM[11799];
assign MEM[36242] = MEM[11696] + MEM[11905];
assign MEM[36243] = MEM[11701] + MEM[12016];
assign MEM[36244] = MEM[11702] + MEM[11710];
assign MEM[36245] = MEM[11706] + MEM[11793];
assign MEM[36246] = MEM[11707] + MEM[12084];
assign MEM[36247] = MEM[11713] + MEM[11837];
assign MEM[36248] = MEM[11716] + MEM[11749];
assign MEM[36249] = MEM[11720] + MEM[11813];
assign MEM[36250] = MEM[11722] + MEM[12029];
assign MEM[36251] = MEM[11724] + MEM[11763];
assign MEM[36252] = MEM[11725] + MEM[11931];
assign MEM[36253] = MEM[11737] + MEM[11787];
assign MEM[36254] = MEM[11740] + MEM[11773];
assign MEM[36255] = MEM[11745] + MEM[11822];
assign MEM[36256] = MEM[11752] + MEM[11791];
assign MEM[36257] = MEM[11754] + MEM[11841];
assign MEM[36258] = MEM[11755] + MEM[11890];
assign MEM[36259] = MEM[11761] + MEM[11830];
assign MEM[36260] = MEM[11766] + MEM[11914];
assign MEM[36261] = MEM[11768] + MEM[11944];
assign MEM[36262] = MEM[11772] + MEM[12223];
assign MEM[36263] = MEM[11778] + MEM[12344];
assign MEM[36264] = MEM[11779] + MEM[11945];
assign MEM[36265] = MEM[11782] + MEM[11854];
assign MEM[36266] = MEM[11784] + MEM[11883];
assign MEM[36267] = MEM[11786] + MEM[11994];
assign MEM[36268] = MEM[11792] + MEM[11933];
assign MEM[36269] = MEM[11800] + MEM[11899];
assign MEM[36270] = MEM[11801] + MEM[12211];
assign MEM[36271] = MEM[11807] + MEM[12152];
assign MEM[36272] = MEM[11808] + MEM[12047];
assign MEM[36273] = MEM[11817] + MEM[11860];
assign MEM[36274] = MEM[11819] + MEM[11861];
assign MEM[36275] = MEM[11826] + MEM[11902];
assign MEM[36276] = MEM[11831] + MEM[12069];
assign MEM[36277] = MEM[11833] + MEM[11838];
assign MEM[36278] = MEM[11834] + MEM[11880];
assign MEM[36279] = MEM[11839] + MEM[11934];
assign MEM[36280] = MEM[11840] + MEM[11865];
assign MEM[36281] = MEM[11847] + MEM[12058];
assign MEM[36282] = MEM[11851] + MEM[11862];
assign MEM[36283] = MEM[11853] + MEM[11892];
assign MEM[36284] = MEM[11856] + MEM[11874];
assign MEM[36285] = MEM[11863] + MEM[12062];
assign MEM[36286] = MEM[11866] + MEM[11967];
assign MEM[36287] = MEM[11868] + MEM[11882];
assign MEM[36288] = MEM[11870] + MEM[11926];
assign MEM[36289] = MEM[11879] + MEM[11885];
assign MEM[36290] = MEM[11888] + MEM[11976];
assign MEM[36291] = MEM[11893] + MEM[11965];
assign MEM[36292] = MEM[11894] + MEM[11922];
assign MEM[36293] = MEM[11896] + MEM[12373];
assign MEM[36294] = MEM[11897] + MEM[11917];
assign MEM[36295] = MEM[11898] + MEM[12079];
assign MEM[36296] = MEM[11907] + MEM[11929];
assign MEM[36297] = MEM[11924] + MEM[12353];
assign MEM[36298] = MEM[11930] + MEM[11940];
assign MEM[36299] = MEM[11932] + MEM[11942];
assign MEM[36300] = MEM[11936] + MEM[12009];
assign MEM[36301] = MEM[11937] + MEM[11943];
assign MEM[36302] = MEM[11939] + MEM[12037];
assign MEM[36303] = MEM[11946] + MEM[11960];
assign MEM[36304] = MEM[11950] + MEM[12355];
assign MEM[36305] = MEM[11954] + MEM[12001];
assign MEM[36306] = MEM[11955] + MEM[11959];
assign MEM[36307] = MEM[11957] + MEM[11958];
assign MEM[36308] = MEM[11961] + MEM[12168];
assign MEM[36309] = MEM[11963] + MEM[12061];
assign MEM[36310] = MEM[11969] + MEM[12191];
assign MEM[36311] = MEM[11972] + MEM[11993];
assign MEM[36312] = MEM[11975] + MEM[11995];
assign MEM[36313] = MEM[11977] + MEM[12013];
assign MEM[36314] = MEM[11978] + MEM[12271];
assign MEM[36315] = MEM[11979] + MEM[11999];
assign MEM[36316] = MEM[11981] + MEM[12039];
assign MEM[36317] = MEM[11985] + MEM[12677];
assign MEM[36318] = MEM[11989] + MEM[12121];
assign MEM[36319] = MEM[11991] + MEM[12025];
assign MEM[36320] = MEM[11992] + MEM[12179];
assign MEM[36321] = MEM[12002] + MEM[12049];
assign MEM[36322] = MEM[12007] + MEM[12349];
assign MEM[36323] = MEM[12010] + MEM[12195];
assign MEM[36324] = MEM[12011] + MEM[12033];
assign MEM[36325] = MEM[12017] + MEM[12160];
assign MEM[36326] = MEM[12019] + MEM[12398];
assign MEM[36327] = MEM[12022] + MEM[12302];
assign MEM[36328] = MEM[12040] + MEM[12138];
assign MEM[36329] = MEM[12046] + MEM[12057];
assign MEM[36330] = MEM[12050] + MEM[12064];
assign MEM[36331] = MEM[12053] + MEM[12374];
assign MEM[36332] = MEM[12059] + MEM[12337];
assign MEM[36333] = MEM[12068] + MEM[12119];
assign MEM[36334] = MEM[12070] + MEM[12454];
assign MEM[36335] = MEM[12073] + MEM[12086];
assign MEM[36336] = MEM[12075] + MEM[12209];
assign MEM[36337] = MEM[12080] + MEM[12200];
assign MEM[36338] = MEM[12087] + MEM[12462];
assign MEM[36339] = MEM[12088] + MEM[12210];
assign MEM[36340] = MEM[12089] + MEM[12128];
assign MEM[36341] = MEM[12091] + MEM[12357];
assign MEM[36342] = MEM[12098] + MEM[12399];
assign MEM[36343] = MEM[12099] + MEM[12851];
assign MEM[36344] = MEM[12104] + MEM[12130];
assign MEM[36345] = MEM[12108] + MEM[12162];
assign MEM[36346] = MEM[12110] + MEM[12149];
assign MEM[36347] = MEM[12113] + MEM[12114];
assign MEM[36348] = MEM[12116] + MEM[12288];
assign MEM[36349] = MEM[12117] + MEM[12247];
assign MEM[36350] = MEM[12126] + MEM[12222];
assign MEM[36351] = MEM[12129] + MEM[12145];
assign MEM[36352] = MEM[12142] + MEM[12285];
assign MEM[36353] = MEM[12144] + MEM[12215];
assign MEM[36354] = MEM[12150] + MEM[12376];
assign MEM[36355] = MEM[12153] + MEM[12331];
assign MEM[36356] = MEM[12154] + MEM[12481];
assign MEM[36357] = MEM[12171] + MEM[12250];
assign MEM[36358] = MEM[12172] + MEM[12369];
assign MEM[36359] = MEM[12180] + MEM[12254];
assign MEM[36360] = MEM[12192] + MEM[12238];
assign MEM[36361] = MEM[12202] + MEM[12445];
assign MEM[36362] = MEM[12213] + MEM[12317];
assign MEM[36363] = MEM[12236] + MEM[12303];
assign MEM[36364] = MEM[12237] + MEM[12408];
assign MEM[36365] = MEM[12240] + MEM[12319];
assign MEM[36366] = MEM[12248] + MEM[12627];
assign MEM[36367] = MEM[12249] + MEM[12397];
assign MEM[36368] = MEM[12260] + MEM[12446];
assign MEM[36369] = MEM[12262] + MEM[12356];
assign MEM[36370] = MEM[12267] + MEM[12368];
assign MEM[36371] = MEM[12269] + MEM[12321];
assign MEM[36372] = MEM[12280] + MEM[12596];
assign MEM[36373] = MEM[12290] + MEM[12527];
assign MEM[36374] = MEM[12295] + MEM[13016];
assign MEM[36375] = MEM[12298] + MEM[12311];
assign MEM[36376] = MEM[12322] + MEM[12613];
assign MEM[36377] = MEM[12336] + MEM[12428];
assign MEM[36378] = MEM[12348] + MEM[12371];
assign MEM[36379] = MEM[12364] + MEM[12402];
assign MEM[36380] = MEM[12365] + MEM[12531];
assign MEM[36381] = MEM[12384] + MEM[12510];
assign MEM[36382] = MEM[12385] + MEM[12453];
assign MEM[36383] = MEM[12389] + MEM[12435];
assign MEM[36384] = MEM[12394] + MEM[12495];
assign MEM[36385] = MEM[12400] + MEM[12617];
assign MEM[36386] = MEM[12401] + MEM[12637];
assign MEM[36387] = MEM[12404] + MEM[12477];
assign MEM[36388] = MEM[12405] + MEM[12571];
assign MEM[36389] = MEM[12410] + MEM[12684];
assign MEM[36390] = MEM[12414] + MEM[12471];
assign MEM[36391] = MEM[12416] + MEM[12452];
assign MEM[36392] = MEM[12420] + MEM[12516];
assign MEM[36393] = MEM[12424] + MEM[12969];
assign MEM[36394] = MEM[12427] + MEM[12482];
assign MEM[36395] = MEM[12430] + MEM[12522];
assign MEM[36396] = MEM[12432] + MEM[12518];
assign MEM[36397] = MEM[12439] + MEM[12680];
assign MEM[36398] = MEM[12440] + MEM[12564];
assign MEM[36399] = MEM[12442] + MEM[12444];
assign MEM[36400] = MEM[12449] + MEM[12548];
assign MEM[36401] = MEM[12450] + MEM[12602];
assign MEM[36402] = MEM[12458] + MEM[12773];
assign MEM[36403] = MEM[12468] + MEM[12493];
assign MEM[36404] = MEM[12475] + MEM[12937];
assign MEM[36405] = MEM[12476] + MEM[12559];
assign MEM[36406] = MEM[12484] + MEM[13132];
assign MEM[36407] = MEM[12485] + MEM[12765];
assign MEM[36408] = MEM[12488] + MEM[12766];
assign MEM[36409] = MEM[12491] + MEM[13104];
assign MEM[36410] = MEM[12505] + MEM[12701];
assign MEM[36411] = MEM[12506] + MEM[12826];
assign MEM[36412] = MEM[12520] + MEM[13114];
assign MEM[36413] = MEM[12521] + MEM[12676];
assign MEM[36414] = MEM[12526] + MEM[12717];
assign MEM[36415] = MEM[12538] + MEM[13442];
assign MEM[36416] = MEM[12541] + MEM[12578];
assign MEM[36417] = MEM[12553] + MEM[13003];
assign MEM[36418] = MEM[12561] + MEM[12752];
assign MEM[36419] = MEM[12567] + MEM[12618];
assign MEM[36420] = MEM[12568] + MEM[12732];
assign MEM[36421] = MEM[12569] + MEM[13054];
assign MEM[36422] = MEM[12574] + MEM[12582];
assign MEM[36423] = MEM[12581] + MEM[12735];
assign MEM[36424] = MEM[12590] + MEM[12768];
assign MEM[36425] = MEM[12592] + MEM[12623];
assign MEM[36426] = MEM[12598] + MEM[12652];
assign MEM[36427] = MEM[12604] + MEM[12829];
assign MEM[36428] = MEM[12611] + MEM[12817];
assign MEM[36429] = MEM[12620] + MEM[12682];
assign MEM[36430] = MEM[12628] + MEM[12747];
assign MEM[36431] = MEM[12631] + MEM[12901];
assign MEM[36432] = MEM[12633] + MEM[12886];
assign MEM[36433] = MEM[12638] + MEM[13215];
assign MEM[36434] = MEM[12649] + MEM[12987];
assign MEM[36435] = MEM[12662] + MEM[12748];
assign MEM[36436] = MEM[12668] + MEM[12921];
assign MEM[36437] = MEM[12672] + MEM[12704];
assign MEM[36438] = MEM[12675] + MEM[12933];
assign MEM[36439] = MEM[12679] + MEM[12688];
assign MEM[36440] = MEM[12681] + MEM[12689];
assign MEM[36441] = MEM[12683] + MEM[12794];
assign MEM[36442] = MEM[12690] + MEM[12938];
assign MEM[36443] = MEM[12693] + MEM[12805];
assign MEM[36444] = MEM[12700] + MEM[12863];
assign MEM[36445] = MEM[12711] + MEM[12720];
assign MEM[36446] = MEM[12715] + MEM[12743];
assign MEM[36447] = MEM[12718] + MEM[13348];
assign MEM[36448] = MEM[12728] + MEM[12842];
assign MEM[36449] = MEM[12729] + MEM[13150];
assign MEM[36450] = MEM[12730] + MEM[12762];
assign MEM[36451] = MEM[12734] + MEM[12860];
assign MEM[36452] = MEM[12756] + MEM[13165];
assign MEM[36453] = MEM[12757] + MEM[12770];
assign MEM[36454] = MEM[12758] + MEM[12819];
assign MEM[36455] = MEM[12763] + MEM[12828];
assign MEM[36456] = MEM[12769] + MEM[13667];
assign MEM[36457] = MEM[12771] + MEM[12979];
assign MEM[36458] = MEM[12781] + MEM[12977];
assign MEM[36459] = MEM[12808] + MEM[13039];
assign MEM[36460] = MEM[12809] + MEM[12838];
assign MEM[36461] = MEM[12812] + MEM[12821];
assign MEM[36462] = MEM[12816] + MEM[13034];
assign MEM[36463] = MEM[12855] + MEM[12945];
assign MEM[36464] = MEM[12865] + MEM[13042];
assign MEM[36465] = MEM[12869] + MEM[12872];
assign MEM[36466] = MEM[12877] + MEM[12918];
assign MEM[36467] = MEM[12878] + MEM[12927];
assign MEM[36468] = MEM[12879] + MEM[13027];
assign MEM[36469] = MEM[12882] + MEM[13199];
assign MEM[36470] = MEM[12887] + MEM[13068];
assign MEM[36471] = MEM[12902] + MEM[12973];
assign MEM[36472] = MEM[12903] + MEM[13072];
assign MEM[36473] = MEM[12905] + MEM[13310];
assign MEM[36474] = MEM[12906] + MEM[12925];
assign MEM[36475] = MEM[12910] + MEM[12950];
assign MEM[36476] = MEM[12911] + MEM[13184];
assign MEM[36477] = MEM[12920] + MEM[13451];
assign MEM[36478] = MEM[12926] + MEM[12994];
assign MEM[36479] = MEM[12928] + MEM[13109];
assign MEM[36480] = MEM[12930] + MEM[13217];
assign MEM[36481] = MEM[12932] + MEM[13007];
assign MEM[36482] = MEM[12947] + MEM[13177];
assign MEM[36483] = MEM[12955] + MEM[13294];
assign MEM[36484] = MEM[12962] + MEM[12972];
assign MEM[36485] = MEM[12963] + MEM[13314];
assign MEM[36486] = MEM[12971] + MEM[13026];
assign MEM[36487] = MEM[12976] + MEM[13062];
assign MEM[36488] = MEM[13001] + MEM[13022];
assign MEM[36489] = MEM[13002] + MEM[13563];
assign MEM[36490] = MEM[13006] + MEM[13409];
assign MEM[36491] = MEM[13008] + MEM[13081];
assign MEM[36492] = MEM[13017] + MEM[13033];
assign MEM[36493] = MEM[13019] + MEM[13164];
assign MEM[36494] = MEM[13025] + MEM[13069];
assign MEM[36495] = MEM[13029] + MEM[13210];
assign MEM[36496] = MEM[13030] + MEM[13558];
assign MEM[36497] = MEM[13032] + MEM[13083];
assign MEM[36498] = MEM[13047] + MEM[13065];
assign MEM[36499] = MEM[13050] + MEM[13098];
assign MEM[36500] = MEM[13052] + MEM[13175];
assign MEM[36501] = MEM[13056] + MEM[13408];
assign MEM[36502] = MEM[13058] + MEM[13102];
assign MEM[36503] = MEM[13061] + MEM[13247];
assign MEM[36504] = MEM[13074] + MEM[13129];
assign MEM[36505] = MEM[13077] + MEM[13136];
assign MEM[36506] = MEM[13084] + MEM[13279];
assign MEM[36507] = MEM[13090] + MEM[13277];
assign MEM[36508] = MEM[13111] + MEM[13204];
assign MEM[36509] = MEM[13125] + MEM[13406];
assign MEM[36510] = MEM[13128] + MEM[13149];
assign MEM[36511] = MEM[13139] + MEM[13671];
assign MEM[36512] = MEM[13140] + MEM[13208];
assign MEM[36513] = MEM[13141] + MEM[13148];
assign MEM[36514] = MEM[13143] + MEM[13392];
assign MEM[36515] = MEM[13154] + MEM[13246];
assign MEM[36516] = MEM[13156] + MEM[13404];
assign MEM[36517] = MEM[13160] + MEM[13313];
assign MEM[36518] = MEM[13176] + MEM[13660];
assign MEM[36519] = MEM[13178] + MEM[13228];
assign MEM[36520] = MEM[13182] + MEM[13231];
assign MEM[36521] = MEM[13193] + MEM[13212];
assign MEM[36522] = MEM[13206] + MEM[13394];
assign MEM[36523] = MEM[13209] + MEM[13317];
assign MEM[36524] = MEM[13221] + MEM[13278];
assign MEM[36525] = MEM[13223] + MEM[13819];
assign MEM[36526] = MEM[13226] + MEM[13367];
assign MEM[36527] = MEM[13227] + MEM[13255];
assign MEM[36528] = MEM[13237] + MEM[13507];
assign MEM[36529] = MEM[13241] + MEM[13252];
assign MEM[36530] = MEM[13244] + MEM[14224];
assign MEM[36531] = MEM[13245] + MEM[13280];
assign MEM[36532] = MEM[13248] + MEM[13287];
assign MEM[36533] = MEM[13256] + MEM[13272];
assign MEM[36534] = MEM[13257] + MEM[13644];
assign MEM[36535] = MEM[13270] + MEM[13293];
assign MEM[36536] = MEM[13271] + MEM[13288];
assign MEM[36537] = MEM[13281] + MEM[13714];
assign MEM[36538] = MEM[13285] + MEM[13436];
assign MEM[36539] = MEM[13290] + MEM[13365];
assign MEM[36540] = MEM[13291] + MEM[13370];
assign MEM[36541] = MEM[13295] + MEM[13301];
assign MEM[36542] = MEM[13300] + MEM[13489];
assign MEM[36543] = MEM[13304] + MEM[13527];
assign MEM[36544] = MEM[13305] + MEM[13397];
assign MEM[36545] = MEM[13307] + MEM[13674];
assign MEM[36546] = MEM[13309] + MEM[13503];
assign MEM[36547] = MEM[13315] + MEM[13391];
assign MEM[36548] = MEM[13330] + MEM[13565];
assign MEM[36549] = MEM[13331] + MEM[13385];
assign MEM[36550] = MEM[13332] + MEM[13333];
assign MEM[36551] = MEM[13335] + MEM[13500];
assign MEM[36552] = MEM[13354] + MEM[13362];
assign MEM[36553] = MEM[13357] + MEM[13461];
assign MEM[36554] = MEM[13363] + MEM[13439];
assign MEM[36555] = MEM[13368] + MEM[13641];
assign MEM[36556] = MEM[13371] + MEM[13381];
assign MEM[36557] = MEM[13373] + MEM[13437];
assign MEM[36558] = MEM[13375] + MEM[13504];
assign MEM[36559] = MEM[13378] + MEM[13589];
assign MEM[36560] = MEM[13387] + MEM[13463];
assign MEM[36561] = MEM[13389] + MEM[13421];
assign MEM[36562] = MEM[13402] + MEM[13441];
assign MEM[36563] = MEM[13416] + MEM[13698];
assign MEM[36564] = MEM[13418] + MEM[13544];
assign MEM[36565] = MEM[13419] + MEM[13426];
assign MEM[36566] = MEM[13422] + MEM[14355];
assign MEM[36567] = MEM[13429] + MEM[13647];
assign MEM[36568] = MEM[13431] + MEM[13576];
assign MEM[36569] = MEM[13434] + MEM[13712];
assign MEM[36570] = MEM[13438] + MEM[13440];
assign MEM[36571] = MEM[13447] + MEM[13499];
assign MEM[36572] = MEM[13453] + MEM[13476];
assign MEM[36573] = MEM[13457] + MEM[13474];
assign MEM[36574] = MEM[13466] + MEM[13724];
assign MEM[36575] = MEM[13469] + MEM[13593];
assign MEM[36576] = MEM[13475] + MEM[13601];
assign MEM[36577] = MEM[13477] + MEM[13478];
assign MEM[36578] = MEM[13480] + MEM[13598];
assign MEM[36579] = MEM[13483] + MEM[13523];
assign MEM[36580] = MEM[13484] + MEM[13596];
assign MEM[36581] = MEM[13492] + MEM[13550];
assign MEM[36582] = MEM[13498] + MEM[13551];
assign MEM[36583] = MEM[13501] + MEM[13640];
assign MEM[36584] = MEM[13502] + MEM[13692];
assign MEM[36585] = MEM[13509] + MEM[13779];
assign MEM[36586] = MEM[13511] + MEM[13619];
assign MEM[36587] = MEM[13518] + MEM[15486];
assign MEM[36588] = MEM[13520] + MEM[15085];
assign MEM[36589] = MEM[13528] + MEM[14023];
assign MEM[36590] = MEM[13533] + MEM[13584];
assign MEM[36591] = MEM[13536] + MEM[14024];
assign MEM[36592] = MEM[13538] + MEM[13887];
assign MEM[36593] = MEM[13547] + MEM[13691];
assign MEM[36594] = MEM[13552] + MEM[13765];
assign MEM[36595] = MEM[13555] + MEM[13747];
assign MEM[36596] = MEM[13556] + MEM[13774];
assign MEM[36597] = MEM[13557] + MEM[15466];
assign MEM[36598] = MEM[13559] + MEM[13574];
assign MEM[36599] = MEM[13560] + MEM[13572];
assign MEM[36600] = MEM[13567] + MEM[13570];
assign MEM[36601] = MEM[13571] + MEM[13679];
assign MEM[36602] = MEM[13575] + MEM[14041];
assign MEM[36603] = MEM[13582] + MEM[13755];
assign MEM[36604] = MEM[13587] + MEM[13811];
assign MEM[36605] = MEM[13592] + MEM[13637];
assign MEM[36606] = MEM[13594] + MEM[13645];
assign MEM[36607] = MEM[13597] + MEM[15583];
assign MEM[36608] = MEM[13599] + MEM[13676];
assign MEM[36609] = MEM[13602] + MEM[13748];
assign MEM[36610] = MEM[13604] + MEM[13695];
assign MEM[36611] = MEM[13606] + MEM[13742];
assign MEM[36612] = MEM[13614] + MEM[13752];
assign MEM[36613] = MEM[13616] + MEM[13706];
assign MEM[36614] = MEM[13621] + MEM[13669];
assign MEM[36615] = MEM[13625] + MEM[13643];
assign MEM[36616] = MEM[13627] + MEM[13713];
assign MEM[36617] = MEM[13628] + MEM[13696];
assign MEM[36618] = MEM[13634] + MEM[15381];
assign MEM[36619] = MEM[13635] + MEM[13678];
assign MEM[36620] = MEM[13639] + MEM[13814];
assign MEM[36621] = MEM[13646] + MEM[15584];
assign MEM[36622] = MEM[13652] + MEM[14263];
assign MEM[36623] = MEM[13655] + MEM[13743];
assign MEM[36624] = MEM[13656] + MEM[13731];
assign MEM[36625] = MEM[13661] + MEM[13708];
assign MEM[36626] = MEM[13668] + MEM[13693];
assign MEM[36627] = MEM[13672] + MEM[13702];
assign MEM[36628] = MEM[13673] + MEM[14278];
assign MEM[36629] = MEM[13682] + MEM[13782];
assign MEM[36630] = MEM[13683] + MEM[13699];
assign MEM[36631] = MEM[13686] + MEM[13727];
assign MEM[36632] = MEM[13689] + MEM[14377];
assign MEM[36633] = MEM[13700] + MEM[13721];
assign MEM[36634] = MEM[13707] + MEM[13973];
assign MEM[36635] = MEM[13710] + MEM[13749];
assign MEM[36636] = MEM[13718] + MEM[13773];
assign MEM[36637] = MEM[13720] + MEM[15272];
assign MEM[36638] = MEM[13722] + MEM[15210];
assign MEM[36639] = MEM[13733] + MEM[13826];
assign MEM[36640] = MEM[13735] + MEM[13839];
assign MEM[36641] = MEM[13737] + MEM[13791];
assign MEM[36642] = MEM[13753] + MEM[14147];
assign MEM[36643] = MEM[13754] + MEM[13849];
assign MEM[36644] = MEM[13756] + MEM[13777];
assign MEM[36645] = MEM[13761] + MEM[13766];
assign MEM[36646] = MEM[13762] + MEM[14771];
assign MEM[36647] = MEM[13764] + MEM[14120];
assign MEM[36648] = MEM[13767] + MEM[14158];
assign MEM[36649] = MEM[13769] + MEM[13770];
assign MEM[36650] = MEM[13775] + MEM[13809];
assign MEM[36651] = MEM[13780] + MEM[13794];
assign MEM[36652] = MEM[13783] + MEM[13963];
assign MEM[36653] = MEM[13785] + MEM[13916];
assign MEM[36654] = MEM[13788] + MEM[15300];
assign MEM[36655] = MEM[13798] + MEM[14008];
assign MEM[36656] = MEM[13799] + MEM[14868];
assign MEM[36657] = MEM[13820] + MEM[13825];
assign MEM[36658] = MEM[13822] + MEM[14384];
assign MEM[36659] = MEM[13823] + MEM[15171];
assign MEM[36660] = MEM[13824] + MEM[14049];
assign MEM[36661] = MEM[13827] + MEM[14310];
assign MEM[36662] = MEM[13897] + MEM[15067];
assign MEM[36663] = MEM[13909] + MEM[14026];
assign MEM[36664] = MEM[13919] + MEM[14221];
assign MEM[36665] = MEM[13939] + MEM[14013];
assign MEM[36666] = MEM[13983] + MEM[15511];
assign MEM[36667] = MEM[13990] + MEM[14559];
assign MEM[36668] = MEM[14009] + MEM[14074];
assign MEM[36669] = MEM[14046] + MEM[14231];
assign MEM[36670] = MEM[14048] + MEM[14079];
assign MEM[36671] = MEM[14078] + MEM[14084];
assign MEM[36672] = MEM[14080] + MEM[14243];
assign MEM[36673] = MEM[14106] + MEM[15671];
assign MEM[36674] = MEM[14117] + MEM[14253];
assign MEM[36675] = MEM[14178] + MEM[14561];
assign MEM[36676] = MEM[14215] + MEM[14641];
assign MEM[36677] = MEM[14217] + MEM[14258];
assign MEM[36678] = MEM[14235] + MEM[14798];
assign MEM[36679] = MEM[14244] + MEM[15611];
assign MEM[36680] = MEM[14273] + MEM[14594];
assign MEM[36681] = MEM[14295] + MEM[15358];
assign MEM[36682] = MEM[14335] + MEM[14389];
assign MEM[36683] = MEM[14387] + MEM[14429];
assign MEM[36684] = MEM[14418] + MEM[14705];
assign MEM[36685] = MEM[14449] + MEM[15701];
assign MEM[36686] = MEM[14464] + MEM[14595];
assign MEM[36687] = MEM[14492] + MEM[14501];
assign MEM[36688] = MEM[14497] + MEM[14966];
assign MEM[36689] = MEM[14517] + MEM[15487];
assign MEM[36690] = MEM[14556] + MEM[15509];
assign MEM[36691] = MEM[14567] + MEM[15385];
assign MEM[36692] = MEM[14575] + MEM[14955];
assign MEM[36693] = MEM[14585] + MEM[14596];
assign MEM[36694] = MEM[14628] + MEM[15710];
assign MEM[36695] = MEM[14630] + MEM[15151];
assign MEM[36696] = MEM[14660] + MEM[15431];
assign MEM[36697] = MEM[14681] + MEM[15080];
assign MEM[36698] = MEM[14691] + MEM[14890];
assign MEM[36699] = MEM[14709] + MEM[15651];
assign MEM[36700] = MEM[14772] + MEM[15563];
assign MEM[36701] = MEM[14784] + MEM[15459];
assign MEM[36702] = MEM[14822] + MEM[15481];
assign MEM[36703] = MEM[14830] + MEM[14928];
assign MEM[36704] = MEM[14871] + MEM[15474];
assign MEM[36705] = MEM[14873] + MEM[14900];
assign MEM[36706] = MEM[14896] + MEM[15025];
assign MEM[36707] = MEM[14902] + MEM[15094];
assign MEM[36708] = MEM[14922] + MEM[15494];
assign MEM[36709] = MEM[14930] + MEM[15184];
assign MEM[36710] = MEM[14992] + MEM[15574];
assign MEM[36711] = MEM[15002] + MEM[15166];
assign MEM[36712] = MEM[15098] + MEM[15211];
assign MEM[36713] = MEM[15100] + MEM[15417];
assign MEM[36714] = MEM[15111] + MEM[15490];
assign MEM[36715] = MEM[15154] + MEM[15538];
assign MEM[36716] = MEM[15163] + MEM[15386];
assign MEM[36717] = MEM[15183] + MEM[15230];
assign MEM[36718] = MEM[15190] + MEM[15332];
assign MEM[36719] = MEM[15191] + MEM[15245];
assign MEM[36720] = MEM[15219] + MEM[15464];
assign MEM[36721] = MEM[15248] + MEM[15361];
assign MEM[36722] = MEM[15270] + MEM[15479];
assign MEM[36723] = MEM[15301] + MEM[15579];
assign MEM[36724] = MEM[15317] + MEM[15626];
assign MEM[36725] = MEM[15330] + MEM[15470];
assign MEM[36726] = MEM[15351] + MEM[15480];
assign MEM[36727] = MEM[15360] + MEM[15427];
assign MEM[36728] = MEM[15374] + MEM[15496];
assign MEM[36729] = MEM[15380] + MEM[15460];
assign MEM[36730] = MEM[15394] + MEM[15695];
assign MEM[36731] = MEM[15403] + MEM[15526];
assign MEM[36732] = MEM[15451] + MEM[15475];
assign MEM[36733] = MEM[15454] + MEM[15468];
assign MEM[36734] = MEM[15456] + MEM[15767];
assign MEM[36735] = MEM[15457] + MEM[15485];
assign MEM[36736] = MEM[15458] + MEM[15737];
assign MEM[36737] = MEM[15462] + MEM[15554];
assign MEM[36738] = MEM[15463] + MEM[15529];
assign MEM[36739] = MEM[15465] + MEM[15540];
assign MEM[36740] = MEM[15467] + MEM[15620];
assign MEM[36741] = MEM[15469] + MEM[15488];
assign MEM[36742] = MEM[15472] + MEM[15683];
assign MEM[36743] = MEM[15476] + MEM[15493];
assign MEM[36744] = MEM[15478] + MEM[15686];
assign MEM[36745] = MEM[15482] + MEM[15539];
assign MEM[36746] = MEM[15483] + MEM[15508];
assign MEM[36747] = MEM[15491] + MEM[15589];
assign MEM[36748] = MEM[15492] + MEM[15499];
assign MEM[36749] = MEM[15497] + MEM[15577];
assign MEM[36750] = MEM[15500] + MEM[15518];
assign MEM[36751] = MEM[15501] + MEM[15569];
assign MEM[36752] = MEM[15505] + MEM[15506];
assign MEM[36753] = MEM[15507] + MEM[15542];
assign MEM[36754] = MEM[15517] + MEM[15536];
assign MEM[36755] = MEM[15519] + MEM[16100];
assign MEM[36756] = MEM[15522] + MEM[15766];
assign MEM[36757] = MEM[15523] + MEM[15730];
assign MEM[36758] = MEM[15524] + MEM[15557];
assign MEM[36759] = MEM[15525] + MEM[15543];
assign MEM[36760] = MEM[15528] + MEM[15772];
assign MEM[36761] = MEM[15530] + MEM[15629];
assign MEM[36762] = MEM[15532] + MEM[15618];
assign MEM[36763] = MEM[15537] + MEM[15650];
assign MEM[36764] = MEM[15545] + MEM[15647];
assign MEM[36765] = MEM[15546] + MEM[15659];
assign MEM[36766] = MEM[15549] + MEM[15564];
assign MEM[36767] = MEM[15550] + MEM[15694];
assign MEM[36768] = MEM[15551] + MEM[15573];
assign MEM[36769] = MEM[15552] + MEM[15677];
assign MEM[36770] = MEM[15553] + MEM[15568];
assign MEM[36771] = MEM[15556] + MEM[15815];
assign MEM[36772] = MEM[15558] + MEM[15608];
assign MEM[36773] = MEM[15559] + MEM[15585];
assign MEM[36774] = MEM[15560] + MEM[15623];
assign MEM[36775] = MEM[15561] + MEM[15648];
assign MEM[36776] = MEM[15565] + MEM[15803];
assign MEM[36777] = MEM[15575] + MEM[15586];
assign MEM[36778] = MEM[15580] + MEM[15752];
assign MEM[36779] = MEM[15581] + MEM[15698];
assign MEM[36780] = MEM[15582] + MEM[15592];
assign MEM[36781] = MEM[15588] + MEM[15704];
assign MEM[36782] = MEM[15593] + MEM[15614];
assign MEM[36783] = MEM[15594] + MEM[15632];
assign MEM[36784] = MEM[15595] + MEM[15846];
assign MEM[36785] = MEM[15597] + MEM[15661];
assign MEM[36786] = MEM[15600] + MEM[15668];
assign MEM[36787] = MEM[15603] + MEM[15954];
assign MEM[36788] = MEM[15604] + MEM[15642];
assign MEM[36789] = MEM[15605] + MEM[15838];
assign MEM[36790] = MEM[15610] + MEM[15681];
assign MEM[36791] = MEM[15613] + MEM[15619];
assign MEM[36792] = MEM[15615] + MEM[15708];
assign MEM[36793] = MEM[15616] + MEM[15697];
assign MEM[36794] = MEM[15621] + MEM[15667];
assign MEM[36795] = MEM[15622] + MEM[15688];
assign MEM[36796] = MEM[15628] + MEM[15711];
assign MEM[36797] = MEM[15630] + MEM[15696];
assign MEM[36798] = MEM[15633] + MEM[15657];
assign MEM[36799] = MEM[15641] + MEM[15768];
assign MEM[36800] = MEM[15643] + MEM[15690];
assign MEM[36801] = MEM[15644] + MEM[15652];
assign MEM[36802] = MEM[15653] + MEM[15655];
assign MEM[36803] = MEM[15654] + MEM[15714];
assign MEM[36804] = MEM[15658] + MEM[15682];
assign MEM[36805] = MEM[15662] + MEM[15736];
assign MEM[36806] = MEM[15669] + MEM[15851];
assign MEM[36807] = MEM[15678] + MEM[15733];
assign MEM[36808] = MEM[15679] + MEM[15727];
assign MEM[36809] = MEM[15685] + MEM[15822];
assign MEM[36810] = MEM[15687] + MEM[15726];
assign MEM[36811] = MEM[15693] + MEM[15712];
assign MEM[36812] = MEM[15699] + MEM[15890];
assign MEM[36813] = MEM[15703] + MEM[15878];
assign MEM[36814] = MEM[15705] + MEM[15748];
assign MEM[36815] = MEM[15706] + MEM[15805];
assign MEM[36816] = MEM[15707] + MEM[15794];
assign MEM[36817] = MEM[15709] + MEM[15734];
assign MEM[36818] = MEM[15718] + MEM[15741];
assign MEM[36819] = MEM[15719] + MEM[15810];
assign MEM[36820] = MEM[15720] + MEM[16002];
assign MEM[36821] = MEM[15721] + MEM[15869];
assign MEM[36822] = MEM[15722] + MEM[15739];
assign MEM[36823] = MEM[15725] + MEM[15970];
assign MEM[36824] = MEM[15728] + MEM[15880];
assign MEM[36825] = MEM[15732] + MEM[15742];
assign MEM[36826] = MEM[15738] + MEM[15777];
assign MEM[36827] = MEM[15740] + MEM[15775];
assign MEM[36828] = MEM[15744] + MEM[15747];
assign MEM[36829] = MEM[15745] + MEM[16022];
assign MEM[36830] = MEM[15751] + MEM[15779];
assign MEM[36831] = MEM[15754] + MEM[16077];
assign MEM[36832] = MEM[15755] + MEM[15758];
assign MEM[36833] = MEM[15757] + MEM[15800];
assign MEM[36834] = MEM[15759] + MEM[15764];
assign MEM[36835] = MEM[15763] + MEM[15806];
assign MEM[36836] = MEM[15765] + MEM[15873];
assign MEM[36837] = MEM[15769] + MEM[16096];
assign MEM[36838] = MEM[15773] + MEM[15782];
assign MEM[36839] = MEM[15781] + MEM[15817];
assign MEM[36840] = MEM[15783] + MEM[15832];
assign MEM[36841] = MEM[15786] + MEM[15879];
assign MEM[36842] = MEM[15789] + MEM[15907];
assign MEM[36843] = MEM[15791] + MEM[15870];
assign MEM[36844] = MEM[15792] + MEM[15839];
assign MEM[36845] = MEM[15795] + MEM[15797];
assign MEM[36846] = MEM[15796] + MEM[15960];
assign MEM[36847] = MEM[15809] + MEM[15858];
assign MEM[36848] = MEM[15811] + MEM[15849];
assign MEM[36849] = MEM[15812] + MEM[15825];
assign MEM[36850] = MEM[15814] + MEM[15885];
assign MEM[36851] = MEM[15818] + MEM[15941];
assign MEM[36852] = MEM[15821] + MEM[15883];
assign MEM[36853] = MEM[15824] + MEM[15840];
assign MEM[36854] = MEM[15828] + MEM[15829];
assign MEM[36855] = MEM[15830] + MEM[15905];
assign MEM[36856] = MEM[15833] + MEM[15874];
assign MEM[36857] = MEM[15834] + MEM[15916];
assign MEM[36858] = MEM[15835] + MEM[15921];
assign MEM[36859] = MEM[15836] + MEM[15850];
assign MEM[36860] = MEM[15837] + MEM[15892];
assign MEM[36861] = MEM[15842] + MEM[16041];
assign MEM[36862] = MEM[15843] + MEM[15855];
assign MEM[36863] = MEM[15854] + MEM[15982];
assign MEM[36864] = MEM[15856] + MEM[15985];
assign MEM[36865] = MEM[15859] + MEM[15950];
assign MEM[36866] = MEM[15862] + MEM[15934];
assign MEM[36867] = MEM[15863] + MEM[15953];
assign MEM[36868] = MEM[15864] + MEM[15887];
assign MEM[36869] = MEM[15866] + MEM[16080];
assign MEM[36870] = MEM[15872] + MEM[15891];
assign MEM[36871] = MEM[15877] + MEM[15901];
assign MEM[36872] = MEM[15881] + MEM[16014];
assign MEM[36873] = MEM[15884] + MEM[15935];
assign MEM[36874] = MEM[15888] + MEM[15981];
assign MEM[36875] = MEM[15889] + MEM[15986];
assign MEM[36876] = MEM[15894] + MEM[15973];
assign MEM[36877] = MEM[15896] + MEM[16042];
assign MEM[36878] = MEM[15898] + MEM[15971];
assign MEM[36879] = MEM[15900] + MEM[16024];
assign MEM[36880] = MEM[15902] + MEM[16016];
assign MEM[36881] = MEM[15904] + MEM[15952];
assign MEM[36882] = MEM[15906] + MEM[16058];
assign MEM[36883] = MEM[15909] + MEM[15955];
assign MEM[36884] = MEM[15911] + MEM[16074];
assign MEM[36885] = MEM[15912] + MEM[15944];
assign MEM[36886] = MEM[15913] + MEM[16027];
assign MEM[36887] = MEM[15915] + MEM[15936];
assign MEM[36888] = MEM[15917] + MEM[15930];
assign MEM[36889] = MEM[15918] + MEM[15988];
assign MEM[36890] = MEM[15919] + MEM[16004];
assign MEM[36891] = MEM[15922] + MEM[16371];
assign MEM[36892] = MEM[15926] + MEM[16068];
assign MEM[36893] = MEM[15928] + MEM[16135];
assign MEM[36894] = MEM[15933] + MEM[16062];
assign MEM[36895] = MEM[15940] + MEM[15959];
assign MEM[36896] = MEM[15943] + MEM[15958];
assign MEM[36897] = MEM[15945] + MEM[15966];
assign MEM[36898] = MEM[15947] + MEM[16153];
assign MEM[36899] = MEM[15949] + MEM[16029];
assign MEM[36900] = MEM[15956] + MEM[15992];
assign MEM[36901] = MEM[15957] + MEM[16115];
assign MEM[36902] = MEM[15961] + MEM[16005];
assign MEM[36903] = MEM[15964] + MEM[16139];
assign MEM[36904] = MEM[15969] + MEM[16015];
assign MEM[36905] = MEM[15972] + MEM[15993];
assign MEM[36906] = MEM[15976] + MEM[15977];
assign MEM[36907] = MEM[15978] + MEM[16930];
assign MEM[36908] = MEM[15979] + MEM[15980];
assign MEM[36909] = MEM[15989] + MEM[16202];
assign MEM[36910] = MEM[15990] + MEM[16012];
assign MEM[36911] = MEM[15991] + MEM[16011];
assign MEM[36912] = MEM[15996] + MEM[16198];
assign MEM[36913] = MEM[15997] + MEM[16076];
assign MEM[36914] = MEM[15998] + MEM[16010];
assign MEM[36915] = MEM[16000] + MEM[16003];
assign MEM[36916] = MEM[16006] + MEM[16048];
assign MEM[36917] = MEM[16017] + MEM[16122];
assign MEM[36918] = MEM[16019] + MEM[16131];
assign MEM[36919] = MEM[16030] + MEM[16304];
assign MEM[36920] = MEM[16032] + MEM[16090];
assign MEM[36921] = MEM[16033] + MEM[16099];
assign MEM[36922] = MEM[16036] + MEM[16053];
assign MEM[36923] = MEM[16037] + MEM[16380];
assign MEM[36924] = MEM[16038] + MEM[16110];
assign MEM[36925] = MEM[16039] + MEM[16167];
assign MEM[36926] = MEM[16043] + MEM[16168];
assign MEM[36927] = MEM[16045] + MEM[16063];
assign MEM[36928] = MEM[16047] + MEM[16254];
assign MEM[36929] = MEM[16050] + MEM[16093];
assign MEM[36930] = MEM[16051] + MEM[16079];
assign MEM[36931] = MEM[16054] + MEM[16186];
assign MEM[36932] = MEM[16055] + MEM[16357];
assign MEM[36933] = MEM[16056] + MEM[16201];
assign MEM[36934] = MEM[16067] + MEM[16101];
assign MEM[36935] = MEM[16069] + MEM[16082];
assign MEM[36936] = MEM[16071] + MEM[16086];
assign MEM[36937] = MEM[16072] + MEM[16092];
assign MEM[36938] = MEM[16075] + MEM[16083];
assign MEM[36939] = MEM[16081] + MEM[16144];
assign MEM[36940] = MEM[16084] + MEM[16174];
assign MEM[36941] = MEM[16088] + MEM[16241];
assign MEM[36942] = MEM[16089] + MEM[16130];
assign MEM[36943] = MEM[16098] + MEM[16105];
assign MEM[36944] = MEM[16106] + MEM[16246];
assign MEM[36945] = MEM[16107] + MEM[16272];
assign MEM[36946] = MEM[16108] + MEM[16111];
assign MEM[36947] = MEM[16109] + MEM[16218];
assign MEM[36948] = MEM[16112] + MEM[16172];
assign MEM[36949] = MEM[16114] + MEM[16154];
assign MEM[36950] = MEM[16116] + MEM[16173];
assign MEM[36951] = MEM[16118] + MEM[16141];
assign MEM[36952] = MEM[16119] + MEM[16320];
assign MEM[36953] = MEM[16120] + MEM[16127];
assign MEM[36954] = MEM[16121] + MEM[16204];
assign MEM[36955] = MEM[16123] + MEM[16455];
assign MEM[36956] = MEM[16124] + MEM[16300];
assign MEM[36957] = MEM[16125] + MEM[16256];
assign MEM[36958] = MEM[16129] + MEM[16251];
assign MEM[36959] = MEM[16132] + MEM[16341];
assign MEM[36960] = MEM[16133] + MEM[16199];
assign MEM[36961] = MEM[16134] + MEM[16288];
assign MEM[36962] = MEM[16136] + MEM[16290];
assign MEM[36963] = MEM[16143] + MEM[16323];
assign MEM[36964] = MEM[16146] + MEM[16208];
assign MEM[36965] = MEM[16148] + MEM[16379];
assign MEM[36966] = MEM[16149] + MEM[16407];
assign MEM[36967] = MEM[16152] + MEM[16639];
assign MEM[36968] = MEM[16155] + MEM[16164];
assign MEM[36969] = MEM[16158] + MEM[16226];
assign MEM[36970] = MEM[16159] + MEM[16298];
assign MEM[36971] = MEM[16161] + MEM[16243];
assign MEM[36972] = MEM[16162] + MEM[16237];
assign MEM[36973] = MEM[16178] + MEM[16216];
assign MEM[36974] = MEM[16179] + MEM[16408];
assign MEM[36975] = MEM[16180] + MEM[16344];
assign MEM[36976] = MEM[16182] + MEM[16220];
assign MEM[36977] = MEM[16184] + MEM[16229];
assign MEM[36978] = MEM[16191] + MEM[16264];
assign MEM[36979] = MEM[16193] + MEM[16370];
assign MEM[36980] = MEM[16205] + MEM[16295];
assign MEM[36981] = MEM[16206] + MEM[16250];
assign MEM[36982] = MEM[16209] + MEM[16410];
assign MEM[36983] = MEM[16210] + MEM[16386];
assign MEM[36984] = MEM[16213] + MEM[16435];
assign MEM[36985] = MEM[16214] + MEM[16384];
assign MEM[36986] = MEM[16219] + MEM[16248];
assign MEM[36987] = MEM[16222] + MEM[16463];
assign MEM[36988] = MEM[16227] + MEM[16271];
assign MEM[36989] = MEM[16230] + MEM[16352];
assign MEM[36990] = MEM[16231] + MEM[16232];
assign MEM[36991] = MEM[16235] + MEM[16378];
assign MEM[36992] = MEM[16236] + MEM[16576];
assign MEM[36993] = MEM[16238] + MEM[16245];
assign MEM[36994] = MEM[16244] + MEM[16343];
assign MEM[36995] = MEM[16260] + MEM[16305];
assign MEM[36996] = MEM[16261] + MEM[16321];
assign MEM[36997] = MEM[16267] + MEM[16281];
assign MEM[36998] = MEM[16269] + MEM[16544];
assign MEM[36999] = MEM[16270] + MEM[16404];
assign MEM[37000] = MEM[16276] + MEM[16347];
assign MEM[37001] = MEM[16278] + MEM[16443];
assign MEM[37002] = MEM[16291] + MEM[16488];
assign MEM[37003] = MEM[16292] + MEM[16429];
assign MEM[37004] = MEM[16294] + MEM[16332];
assign MEM[37005] = MEM[16297] + MEM[16306];
assign MEM[37006] = MEM[16299] + MEM[16336];
assign MEM[37007] = MEM[16303] + MEM[16467];
assign MEM[37008] = MEM[16308] + MEM[16312];
assign MEM[37009] = MEM[16310] + MEM[16349];
assign MEM[37010] = MEM[16311] + MEM[16568];
assign MEM[37011] = MEM[16313] + MEM[16356];
assign MEM[37012] = MEM[16314] + MEM[16333];
assign MEM[37013] = MEM[16315] + MEM[16330];
assign MEM[37014] = MEM[16318] + MEM[16322];
assign MEM[37015] = MEM[16319] + MEM[16359];
assign MEM[37016] = MEM[16325] + MEM[16360];
assign MEM[37017] = MEM[16327] + MEM[16417];
assign MEM[37018] = MEM[16328] + MEM[16598];
assign MEM[37019] = MEM[16329] + MEM[16556];
assign MEM[37020] = MEM[16331] + MEM[16474];
assign MEM[37021] = MEM[16337] + MEM[16346];
assign MEM[37022] = MEM[16345] + MEM[16382];
assign MEM[37023] = MEM[16348] + MEM[16594];
assign MEM[37024] = MEM[16350] + MEM[16365];
assign MEM[37025] = MEM[16351] + MEM[16374];
assign MEM[37026] = MEM[16353] + MEM[16362];
assign MEM[37027] = MEM[16361] + MEM[16412];
assign MEM[37028] = MEM[16372] + MEM[16444];
assign MEM[37029] = MEM[16373] + MEM[16385];
assign MEM[37030] = MEM[16375] + MEM[16449];
assign MEM[37031] = MEM[16383] + MEM[16477];
assign MEM[37032] = MEM[16387] + MEM[16459];
assign MEM[37033] = MEM[16391] + MEM[16451];
assign MEM[37034] = MEM[16392] + MEM[16581];
assign MEM[37035] = MEM[16395] + MEM[16465];
assign MEM[37036] = MEM[16396] + MEM[16648];
assign MEM[37037] = MEM[16398] + MEM[16454];
assign MEM[37038] = MEM[16399] + MEM[16507];
assign MEM[37039] = MEM[16405] + MEM[16447];
assign MEM[37040] = MEM[16406] + MEM[16428];
assign MEM[37041] = MEM[16409] + MEM[16458];
assign MEM[37042] = MEM[16413] + MEM[16461];
assign MEM[37043] = MEM[16415] + MEM[16416];
assign MEM[37044] = MEM[16419] + MEM[16528];
assign MEM[37045] = MEM[16421] + MEM[16557];
assign MEM[37046] = MEM[16426] + MEM[16710];
assign MEM[37047] = MEM[16430] + MEM[16453];
assign MEM[37048] = MEM[16431] + MEM[16554];
assign MEM[37049] = MEM[16433] + MEM[16622];
assign MEM[37050] = MEM[16437] + MEM[16530];
assign MEM[37051] = MEM[16440] + MEM[16487];
assign MEM[37052] = MEM[16441] + MEM[16608];
assign MEM[37053] = MEM[16445] + MEM[16586];
assign MEM[37054] = MEM[16457] + MEM[16466];
assign MEM[37055] = MEM[16462] + MEM[16607];
assign MEM[37056] = MEM[16464] + MEM[16486];
assign MEM[37057] = MEM[16468] + MEM[16596];
assign MEM[37058] = MEM[16469] + MEM[16490];
assign MEM[37059] = MEM[16471] + MEM[16475];
assign MEM[37060] = MEM[16472] + MEM[16687];
assign MEM[37061] = MEM[16473] + MEM[16663];
assign MEM[37062] = MEM[16476] + MEM[16523];
assign MEM[37063] = MEM[16479] + MEM[16714];
assign MEM[37064] = MEM[16480] + MEM[16712];
assign MEM[37065] = MEM[16482] + MEM[16584];
assign MEM[37066] = MEM[16485] + MEM[16492];
assign MEM[37067] = MEM[16489] + MEM[16506];
assign MEM[37068] = MEM[16491] + MEM[16540];
assign MEM[37069] = MEM[16494] + MEM[16512];
assign MEM[37070] = MEM[16495] + MEM[16906];
assign MEM[37071] = MEM[16496] + MEM[16696];
assign MEM[37072] = MEM[16497] + MEM[16529];
assign MEM[37073] = MEM[16498] + MEM[16570];
assign MEM[37074] = MEM[16503] + MEM[16623];
assign MEM[37075] = MEM[16505] + MEM[16558];
assign MEM[37076] = MEM[16508] + MEM[16519];
assign MEM[37077] = MEM[16511] + MEM[16537];
assign MEM[37078] = MEM[16515] + MEM[16617];
assign MEM[37079] = MEM[16522] + MEM[16572];
assign MEM[37080] = MEM[16524] + MEM[16592];
assign MEM[37081] = MEM[16543] + MEM[16582];
assign MEM[37082] = MEM[16545] + MEM[16580];
assign MEM[37083] = MEM[16550] + MEM[16604];
assign MEM[37084] = MEM[16553] + MEM[16655];
assign MEM[37085] = MEM[16559] + MEM[16635];
assign MEM[37086] = MEM[16564] + MEM[16643];
assign MEM[37087] = MEM[16567] + MEM[16882];
assign MEM[37088] = MEM[16574] + MEM[16590];
assign MEM[37089] = MEM[16578] + MEM[16664];
assign MEM[37090] = MEM[16583] + MEM[16616];
assign MEM[37091] = MEM[16589] + MEM[16727];
assign MEM[37092] = MEM[16591] + MEM[16613];
assign MEM[37093] = MEM[16593] + MEM[16597];
assign MEM[37094] = MEM[16599] + MEM[16699];
assign MEM[37095] = MEM[16601] + MEM[16905];
assign MEM[37096] = MEM[16609] + MEM[16978];
assign MEM[37097] = MEM[16610] + MEM[16659];
assign MEM[37098] = MEM[16615] + MEM[16726];
assign MEM[37099] = MEM[16618] + MEM[16721];
assign MEM[37100] = MEM[16619] + MEM[16637];
assign MEM[37101] = MEM[16625] + MEM[16626];
assign MEM[37102] = MEM[16629] + MEM[16707];
assign MEM[37103] = MEM[16631] + MEM[16677];
assign MEM[37104] = MEM[16633] + MEM[16716];
assign MEM[37105] = MEM[16641] + MEM[16649];
assign MEM[37106] = MEM[16642] + MEM[16653];
assign MEM[37107] = MEM[16646] + MEM[16937];
assign MEM[37108] = MEM[16647] + MEM[16666];
assign MEM[37109] = MEM[16652] + MEM[16792];
assign MEM[37110] = MEM[16658] + MEM[16671];
assign MEM[37111] = MEM[16660] + MEM[16684];
assign MEM[37112] = MEM[16661] + MEM[16680];
assign MEM[37113] = MEM[16667] + MEM[16761];
assign MEM[37114] = MEM[16668] + MEM[17230];
assign MEM[37115] = MEM[16669] + MEM[16679];
assign MEM[37116] = MEM[16672] + MEM[16801];
assign MEM[37117] = MEM[16673] + MEM[16802];
assign MEM[37118] = MEM[16674] + MEM[16749];
assign MEM[37119] = MEM[16675] + MEM[16676];
assign MEM[37120] = MEM[16678] + MEM[17077];
assign MEM[37121] = MEM[16681] + MEM[16715];
assign MEM[37122] = MEM[16682] + MEM[16772];
assign MEM[37123] = MEM[16688] + MEM[16706];
assign MEM[37124] = MEM[16689] + MEM[16690];
assign MEM[37125] = MEM[16692] + MEM[16817];
assign MEM[37126] = MEM[16693] + MEM[16782];
assign MEM[37127] = MEM[16697] + MEM[16732];
assign MEM[37128] = MEM[16698] + MEM[16724];
assign MEM[37129] = MEM[16705] + MEM[16708];
assign MEM[37130] = MEM[16709] + MEM[17110];
assign MEM[37131] = MEM[16713] + MEM[16975];
assign MEM[37132] = MEM[16717] + MEM[16719];
assign MEM[37133] = MEM[16720] + MEM[16805];
assign MEM[37134] = MEM[16722] + MEM[16824];
assign MEM[37135] = MEM[16725] + MEM[16816];
assign MEM[37136] = MEM[16728] + MEM[16773];
assign MEM[37137] = MEM[16729] + MEM[16885];
assign MEM[37138] = MEM[16730] + MEM[16751];
assign MEM[37139] = MEM[16735] + MEM[16837];
assign MEM[37140] = MEM[16737] + MEM[16756];
assign MEM[37141] = MEM[16742] + MEM[16951];
assign MEM[37142] = MEM[16744] + MEM[16858];
assign MEM[37143] = MEM[16745] + MEM[16826];
assign MEM[37144] = MEM[16747] + MEM[16755];
assign MEM[37145] = MEM[16748] + MEM[16758];
assign MEM[37146] = MEM[16753] + MEM[16775];
assign MEM[37147] = MEM[16757] + MEM[16811];
assign MEM[37148] = MEM[16763] + MEM[16812];
assign MEM[37149] = MEM[16765] + MEM[16903];
assign MEM[37150] = MEM[16766] + MEM[17112];
assign MEM[37151] = MEM[16770] + MEM[16793];
assign MEM[37152] = MEM[16771] + MEM[16907];
assign MEM[37153] = MEM[16774] + MEM[17251];
assign MEM[37154] = MEM[16776] + MEM[17182];
assign MEM[37155] = MEM[16781] + MEM[16942];
assign MEM[37156] = MEM[16789] + MEM[16832];
assign MEM[37157] = MEM[16794] + MEM[16898];
assign MEM[37158] = MEM[16797] + MEM[16941];
assign MEM[37159] = MEM[16799] + MEM[16814];
assign MEM[37160] = MEM[16800] + MEM[16895];
assign MEM[37161] = MEM[16803] + MEM[16815];
assign MEM[37162] = MEM[16804] + MEM[17095];
assign MEM[37163] = MEM[16806] + MEM[16852];
assign MEM[37164] = MEM[16810] + MEM[16859];
assign MEM[37165] = MEM[16819] + MEM[16827];
assign MEM[37166] = MEM[16820] + MEM[16828];
assign MEM[37167] = MEM[16822] + MEM[16851];
assign MEM[37168] = MEM[16829] + MEM[16901];
assign MEM[37169] = MEM[16830] + MEM[17119];
assign MEM[37170] = MEM[16834] + MEM[16845];
assign MEM[37171] = MEM[16835] + MEM[16874];
assign MEM[37172] = MEM[16841] + MEM[16925];
assign MEM[37173] = MEM[16842] + MEM[16929];
assign MEM[37174] = MEM[16843] + MEM[17010];
assign MEM[37175] = MEM[16844] + MEM[16883];
assign MEM[37176] = MEM[16849] + MEM[16880];
assign MEM[37177] = MEM[16853] + MEM[16921];
assign MEM[37178] = MEM[16854] + MEM[16936];
assign MEM[37179] = MEM[16855] + MEM[17034];
assign MEM[37180] = MEM[16861] + MEM[16909];
assign MEM[37181] = MEM[16862] + MEM[16923];
assign MEM[37182] = MEM[16869] + MEM[16946];
assign MEM[37183] = MEM[16870] + MEM[16971];
assign MEM[37184] = MEM[16871] + MEM[16889];
assign MEM[37185] = MEM[16873] + MEM[16919];
assign MEM[37186] = MEM[16877] + MEM[16886];
assign MEM[37187] = MEM[16881] + MEM[16893];
assign MEM[37188] = MEM[16887] + MEM[16966];
assign MEM[37189] = MEM[16888] + MEM[16920];
assign MEM[37190] = MEM[16890] + MEM[16913];
assign MEM[37191] = MEM[16896] + MEM[17192];
assign MEM[37192] = MEM[16897] + MEM[16950];
assign MEM[37193] = MEM[16899] + MEM[17000];
assign MEM[37194] = MEM[16900] + MEM[16969];
assign MEM[37195] = MEM[16910] + MEM[17023];
assign MEM[37196] = MEM[16922] + MEM[17199];
assign MEM[37197] = MEM[16924] + MEM[16938];
assign MEM[37198] = MEM[16928] + MEM[17331];
assign MEM[37199] = MEM[16931] + MEM[17103];
assign MEM[37200] = MEM[16933] + MEM[16990];
assign MEM[37201] = MEM[16934] + MEM[17016];
assign MEM[37202] = MEM[16940] + MEM[17144];
assign MEM[37203] = MEM[16944] + MEM[17049];
assign MEM[37204] = MEM[16945] + MEM[17022];
assign MEM[37205] = MEM[16947] + MEM[17108];
assign MEM[37206] = MEM[16948] + MEM[17116];
assign MEM[37207] = MEM[16949] + MEM[16986];
assign MEM[37208] = MEM[16960] + MEM[16979];
assign MEM[37209] = MEM[16964] + MEM[16995];
assign MEM[37210] = MEM[16965] + MEM[17026];
assign MEM[37211] = MEM[16970] + MEM[16992];
assign MEM[37212] = MEM[16972] + MEM[17155];
assign MEM[37213] = MEM[16973] + MEM[17139];
assign MEM[37214] = MEM[16974] + MEM[17018];
assign MEM[37215] = MEM[16976] + MEM[17389];
assign MEM[37216] = MEM[16977] + MEM[17021];
assign MEM[37217] = MEM[16980] + MEM[17042];
assign MEM[37218] = MEM[16981] + MEM[17089];
assign MEM[37219] = MEM[16982] + MEM[17117];
assign MEM[37220] = MEM[16983] + MEM[17140];
assign MEM[37221] = MEM[16984] + MEM[17156];
assign MEM[37222] = MEM[16988] + MEM[17515];
assign MEM[37223] = MEM[16991] + MEM[17048];
assign MEM[37224] = MEM[16993] + MEM[17059];
assign MEM[37225] = MEM[16998] + MEM[17012];
assign MEM[37226] = MEM[17001] + MEM[17037];
assign MEM[37227] = MEM[17004] + MEM[17191];
assign MEM[37228] = MEM[17005] + MEM[17250];
assign MEM[37229] = MEM[17008] + MEM[17027];
assign MEM[37230] = MEM[17011] + MEM[17043];
assign MEM[37231] = MEM[17015] + MEM[17189];
assign MEM[37232] = MEM[17025] + MEM[17130];
assign MEM[37233] = MEM[17030] + MEM[17221];
assign MEM[37234] = MEM[17031] + MEM[17444];
assign MEM[37235] = MEM[17036] + MEM[17127];
assign MEM[37236] = MEM[17039] + MEM[17162];
assign MEM[37237] = MEM[17040] + MEM[17167];
assign MEM[37238] = MEM[17044] + MEM[17128];
assign MEM[37239] = MEM[17047] + MEM[17163];
assign MEM[37240] = MEM[17055] + MEM[17087];
assign MEM[37241] = MEM[17057] + MEM[17066];
assign MEM[37242] = MEM[17060] + MEM[17079];
assign MEM[37243] = MEM[17062] + MEM[17194];
assign MEM[37244] = MEM[17064] + MEM[17455];
assign MEM[37245] = MEM[17069] + MEM[17142];
assign MEM[37246] = MEM[17070] + MEM[17248];
assign MEM[37247] = MEM[17071] + MEM[17076];
assign MEM[37248] = MEM[17073] + MEM[17081];
assign MEM[37249] = MEM[17074] + MEM[17457];
assign MEM[37250] = MEM[17078] + MEM[17366];
assign MEM[37251] = MEM[17086] + MEM[17217];
assign MEM[37252] = MEM[17091] + MEM[17135];
assign MEM[37253] = MEM[17094] + MEM[17242];
assign MEM[37254] = MEM[17098] + MEM[17346];
assign MEM[37255] = MEM[17100] + MEM[17178];
assign MEM[37256] = MEM[17105] + MEM[17241];
assign MEM[37257] = MEM[17106] + MEM[17414];
assign MEM[37258] = MEM[17107] + MEM[17359];
assign MEM[37259] = MEM[17109] + MEM[17157];
assign MEM[37260] = MEM[17111] + MEM[17188];
assign MEM[37261] = MEM[17114] + MEM[17141];
assign MEM[37262] = MEM[17120] + MEM[17129];
assign MEM[37263] = MEM[17124] + MEM[17362];
assign MEM[37264] = MEM[17126] + MEM[17497];
assign MEM[37265] = MEM[17131] + MEM[17138];
assign MEM[37266] = MEM[17137] + MEM[17243];
assign MEM[37267] = MEM[17145] + MEM[17186];
assign MEM[37268] = MEM[17148] + MEM[17271];
assign MEM[37269] = MEM[17151] + MEM[17177];
assign MEM[37270] = MEM[17158] + MEM[17172];
assign MEM[37271] = MEM[17159] + MEM[17256];
assign MEM[37272] = MEM[17160] + MEM[17164];
assign MEM[37273] = MEM[17161] + MEM[17236];
assign MEM[37274] = MEM[17165] + MEM[17293];
assign MEM[37275] = MEM[17168] + MEM[17220];
assign MEM[37276] = MEM[17174] + MEM[17321];
assign MEM[37277] = MEM[17175] + MEM[17336];
assign MEM[37278] = MEM[17184] + MEM[17289];
assign MEM[37279] = MEM[17193] + MEM[17228];
assign MEM[37280] = MEM[17195] + MEM[17388];
assign MEM[37281] = MEM[17196] + MEM[17235];
assign MEM[37282] = MEM[17204] + MEM[17316];
assign MEM[37283] = MEM[17206] + MEM[17232];
assign MEM[37284] = MEM[17208] + MEM[17240];
assign MEM[37285] = MEM[17210] + MEM[17249];
assign MEM[37286] = MEM[17213] + MEM[17258];
assign MEM[37287] = MEM[17215] + MEM[17268];
assign MEM[37288] = MEM[17216] + MEM[17498];
assign MEM[37289] = MEM[17219] + MEM[17501];
assign MEM[37290] = MEM[17223] + MEM[17247];
assign MEM[37291] = MEM[17224] + MEM[17254];
assign MEM[37292] = MEM[17225] + MEM[17303];
assign MEM[37293] = MEM[17226] + MEM[17285];
assign MEM[37294] = MEM[17229] + MEM[17506];
assign MEM[37295] = MEM[17233] + MEM[17253];
assign MEM[37296] = MEM[17234] + MEM[17342];
assign MEM[37297] = MEM[17244] + MEM[17399];
assign MEM[37298] = MEM[17252] + MEM[17560];
assign MEM[37299] = MEM[17255] + MEM[17340];
assign MEM[37300] = MEM[17259] + MEM[17350];
assign MEM[37301] = MEM[17261] + MEM[17479];
assign MEM[37302] = MEM[17265] + MEM[17343];
assign MEM[37303] = MEM[17270] + MEM[17426];
assign MEM[37304] = MEM[17274] + MEM[17281];
assign MEM[37305] = MEM[17275] + MEM[17355];
assign MEM[37306] = MEM[17276] + MEM[17287];
assign MEM[37307] = MEM[17277] + MEM[17341];
assign MEM[37308] = MEM[17278] + MEM[17288];
assign MEM[37309] = MEM[17283] + MEM[17324];
assign MEM[37310] = MEM[17291] + MEM[17351];
assign MEM[37311] = MEM[17295] + MEM[17580];
assign MEM[37312] = MEM[17299] + MEM[17587];
assign MEM[37313] = MEM[17300] + MEM[17301];
assign MEM[37314] = MEM[17302] + MEM[17433];
assign MEM[37315] = MEM[17306] + MEM[17443];
assign MEM[37316] = MEM[17309] + MEM[17360];
assign MEM[37317] = MEM[17311] + MEM[17380];
assign MEM[37318] = MEM[17314] + MEM[17337];
assign MEM[37319] = MEM[17317] + MEM[17448];
assign MEM[37320] = MEM[17320] + MEM[17459];
assign MEM[37321] = MEM[17327] + MEM[17392];
assign MEM[37322] = MEM[17335] + MEM[17517];
assign MEM[37323] = MEM[17344] + MEM[17449];
assign MEM[37324] = MEM[17345] + MEM[17361];
assign MEM[37325] = MEM[17347] + MEM[17484];
assign MEM[37326] = MEM[17348] + MEM[17458];
assign MEM[37327] = MEM[17357] + MEM[17409];
assign MEM[37328] = MEM[17363] + MEM[17746];
assign MEM[37329] = MEM[17367] + MEM[17391];
assign MEM[37330] = MEM[17371] + MEM[17386];
assign MEM[37331] = MEM[17372] + MEM[17375];
assign MEM[37332] = MEM[17374] + MEM[17397];
assign MEM[37333] = MEM[17377] + MEM[17390];
assign MEM[37334] = MEM[17381] + MEM[17503];
assign MEM[37335] = MEM[17384] + MEM[17480];
assign MEM[37336] = MEM[17393] + MEM[17702];
assign MEM[37337] = MEM[17394] + MEM[17593];
assign MEM[37338] = MEM[17395] + MEM[17471];
assign MEM[37339] = MEM[17396] + MEM[17476];
assign MEM[37340] = MEM[17400] + MEM[17541];
assign MEM[37341] = MEM[17408] + MEM[17653];
assign MEM[37342] = MEM[17410] + MEM[17431];
assign MEM[37343] = MEM[17413] + MEM[17703];
assign MEM[37344] = MEM[17415] + MEM[17530];
assign MEM[37345] = MEM[17418] + MEM[17421];
assign MEM[37346] = MEM[17420] + MEM[17516];
assign MEM[37347] = MEM[17425] + MEM[17435];
assign MEM[37348] = MEM[17437] + MEM[17493];
assign MEM[37349] = MEM[17450] + MEM[17451];
assign MEM[37350] = MEM[17453] + MEM[17491];
assign MEM[37351] = MEM[17454] + MEM[17527];
assign MEM[37352] = MEM[17462] + MEM[17495];
assign MEM[37353] = MEM[17464] + MEM[17673];
assign MEM[37354] = MEM[17468] + MEM[17469];
assign MEM[37355] = MEM[17472] + MEM[17483];
assign MEM[37356] = MEM[17477] + MEM[17688];
assign MEM[37357] = MEM[17478] + MEM[17511];
assign MEM[37358] = MEM[17481] + MEM[17509];
assign MEM[37359] = MEM[17486] + MEM[17502];
assign MEM[37360] = MEM[17487] + MEM[17522];
assign MEM[37361] = MEM[17489] + MEM[17510];
assign MEM[37362] = MEM[17490] + MEM[17568];
assign MEM[37363] = MEM[17492] + MEM[17521];
assign MEM[37364] = MEM[17494] + MEM[17520];
assign MEM[37365] = MEM[17496] + MEM[17546];
assign MEM[37366] = MEM[17499] + MEM[17631];
assign MEM[37367] = MEM[17500] + MEM[17538];
assign MEM[37368] = MEM[17504] + MEM[17596];
assign MEM[37369] = MEM[17505] + MEM[17583];
assign MEM[37370] = MEM[17507] + MEM[17551];
assign MEM[37371] = MEM[17508] + MEM[17615];
assign MEM[37372] = MEM[17512] + MEM[17561];
assign MEM[37373] = MEM[17513] + MEM[17526];
assign MEM[37374] = MEM[17514] + MEM[17571];
assign MEM[37375] = MEM[17518] + MEM[17549];
assign MEM[37376] = MEM[17519] + MEM[17575];
assign MEM[37377] = MEM[17523] + MEM[17533];
assign MEM[37378] = MEM[17524] + MEM[17701];
assign MEM[37379] = MEM[17525] + MEM[17655];
assign MEM[37380] = MEM[17528] + MEM[17718];
assign MEM[37381] = MEM[17531] + MEM[17566];
assign MEM[37382] = MEM[17536] + MEM[17687];
assign MEM[37383] = MEM[17537] + MEM[17574];
assign MEM[37384] = MEM[17540] + MEM[17611];
assign MEM[37385] = MEM[17542] + MEM[17544];
assign MEM[37386] = MEM[17543] + MEM[17586];
assign MEM[37387] = MEM[17545] + MEM[17626];
assign MEM[37388] = MEM[17547] + MEM[17592];
assign MEM[37389] = MEM[17548] + MEM[17572];
assign MEM[37390] = MEM[17550] + MEM[17597];
assign MEM[37391] = MEM[17552] + MEM[17676];
assign MEM[37392] = MEM[17553] + MEM[17624];
assign MEM[37393] = MEM[17554] + MEM[17774];
assign MEM[37394] = MEM[17555] + MEM[17569];
assign MEM[37395] = MEM[17557] + MEM[17558];
assign MEM[37396] = MEM[17562] + MEM[17612];
assign MEM[37397] = MEM[17564] + MEM[17753];
assign MEM[37398] = MEM[17570] + MEM[17720];
assign MEM[37399] = MEM[17577] + MEM[17610];
assign MEM[37400] = MEM[17578] + MEM[17671];
assign MEM[37401] = MEM[17579] + MEM[17632];
assign MEM[37402] = MEM[17581] + MEM[17620];
assign MEM[37403] = MEM[17582] + MEM[17649];
assign MEM[37404] = MEM[17584] + MEM[17617];
assign MEM[37405] = MEM[17588] + MEM[17591];
assign MEM[37406] = MEM[17589] + MEM[17694];
assign MEM[37407] = MEM[17590] + MEM[17686];
assign MEM[37408] = MEM[17594] + MEM[17712];
assign MEM[37409] = MEM[17595] + MEM[17599];
assign MEM[37410] = MEM[17598] + MEM[17663];
assign MEM[37411] = MEM[17601] + MEM[17797];
assign MEM[37412] = MEM[17603] + MEM[17656];
assign MEM[37413] = MEM[17604] + MEM[17640];
assign MEM[37414] = MEM[17605] + MEM[17635];
assign MEM[37415] = MEM[17606] + MEM[17634];
assign MEM[37416] = MEM[17607] + MEM[17613];
assign MEM[37417] = MEM[17608] + MEM[17616];
assign MEM[37418] = MEM[17609] + MEM[17817];
assign MEM[37419] = MEM[17614] + MEM[17651];
assign MEM[37420] = MEM[17618] + MEM[17622];
assign MEM[37421] = MEM[17619] + MEM[17737];
assign MEM[37422] = MEM[17621] + MEM[17630];
assign MEM[37423] = MEM[17628] + MEM[17724];
assign MEM[37424] = MEM[17633] + MEM[17762];
assign MEM[37425] = MEM[17636] + MEM[17646];
assign MEM[37426] = MEM[17637] + MEM[17744];
assign MEM[37427] = MEM[17638] + MEM[17652];
assign MEM[37428] = MEM[17639] + MEM[17648];
assign MEM[37429] = MEM[17641] + MEM[17705];
assign MEM[37430] = MEM[17642] + MEM[17665];
assign MEM[37431] = MEM[17643] + MEM[17661];
assign MEM[37432] = MEM[17644] + MEM[17669];
assign MEM[37433] = MEM[17647] + MEM[17689];
assign MEM[37434] = MEM[17650] + MEM[17721];
assign MEM[37435] = MEM[17654] + MEM[17677];
assign MEM[37436] = MEM[17657] + MEM[17698];
assign MEM[37437] = MEM[17658] + MEM[17997];
assign MEM[37438] = MEM[17659] + MEM[17771];
assign MEM[37439] = MEM[17660] + MEM[17691];
assign MEM[37440] = MEM[17664] + MEM[17674];
assign MEM[37441] = MEM[17668] + MEM[17681];
assign MEM[37442] = MEM[17670] + MEM[17760];
assign MEM[37443] = MEM[17675] + MEM[17815];
assign MEM[37444] = MEM[17678] + MEM[17683];
assign MEM[37445] = MEM[17679] + MEM[17697];
assign MEM[37446] = MEM[17680] + MEM[17809];
assign MEM[37447] = MEM[17682] + MEM[17776];
assign MEM[37448] = MEM[17684] + MEM[17854];
assign MEM[37449] = MEM[17685] + MEM[17790];
assign MEM[37450] = MEM[17690] + MEM[17826];
assign MEM[37451] = MEM[17692] + MEM[17779];
assign MEM[37452] = MEM[17699] + MEM[17775];
assign MEM[37453] = MEM[17700] + MEM[17745];
assign MEM[37454] = MEM[17704] + MEM[17766];
assign MEM[37455] = MEM[17706] + MEM[17838];
assign MEM[37456] = MEM[17708] + MEM[17770];
assign MEM[37457] = MEM[17711] + MEM[17748];
assign MEM[37458] = MEM[17714] + MEM[17727];
assign MEM[37459] = MEM[17715] + MEM[17890];
assign MEM[37460] = MEM[17717] + MEM[17788];
assign MEM[37461] = MEM[17719] + MEM[17749];
assign MEM[37462] = MEM[17722] + MEM[17836];
assign MEM[37463] = MEM[17725] + MEM[17785];
assign MEM[37464] = MEM[17726] + MEM[17803];
assign MEM[37465] = MEM[17728] + MEM[17738];
assign MEM[37466] = MEM[17729] + MEM[17840];
assign MEM[37467] = MEM[17730] + MEM[17862];
assign MEM[37468] = MEM[17733] + MEM[17805];
assign MEM[37469] = MEM[17735] + MEM[17763];
assign MEM[37470] = MEM[17736] + MEM[17846];
assign MEM[37471] = MEM[17739] + MEM[17954];
assign MEM[37472] = MEM[17741] + MEM[17828];
assign MEM[37473] = MEM[17743] + MEM[17755];
assign MEM[37474] = MEM[17750] + MEM[17767];
assign MEM[37475] = MEM[17751] + MEM[17849];
assign MEM[37476] = MEM[17752] + MEM[17764];
assign MEM[37477] = MEM[17761] + MEM[17792];
assign MEM[37478] = MEM[17765] + MEM[17780];
assign MEM[37479] = MEM[17768] + MEM[17931];
assign MEM[37480] = MEM[17772] + MEM[17969];
assign MEM[37481] = MEM[17773] + MEM[17798];
assign MEM[37482] = MEM[17777] + MEM[17793];
assign MEM[37483] = MEM[17778] + MEM[17834];
assign MEM[37484] = MEM[17781] + MEM[17787];
assign MEM[37485] = MEM[17783] + MEM[17855];
assign MEM[37486] = MEM[17784] + MEM[17874];
assign MEM[37487] = MEM[17789] + MEM[17830];
assign MEM[37488] = MEM[17791] + MEM[17909];
assign MEM[37489] = MEM[17794] + MEM[17816];
assign MEM[37490] = MEM[17795] + MEM[17821];
assign MEM[37491] = MEM[17800] + MEM[17825];
assign MEM[37492] = MEM[17801] + MEM[17938];
assign MEM[37493] = MEM[17802] + MEM[17875];
assign MEM[37494] = MEM[17804] + MEM[17810];
assign MEM[37495] = MEM[17807] + MEM[17960];
assign MEM[37496] = MEM[17811] + MEM[17843];
assign MEM[37497] = MEM[17812] + MEM[17882];
assign MEM[37498] = MEM[17814] + MEM[17913];
assign MEM[37499] = MEM[17818] + MEM[18110];
assign MEM[37500] = MEM[17819] + MEM[17859];
assign MEM[37501] = MEM[17820] + MEM[17848];
assign MEM[37502] = MEM[17823] + MEM[17873];
assign MEM[37503] = MEM[17824] + MEM[17860];
assign MEM[37504] = MEM[17829] + MEM[17991];
assign MEM[37505] = MEM[17831] + MEM[17892];
assign MEM[37506] = MEM[17833] + MEM[17835];
assign MEM[37507] = MEM[17837] + MEM[17948];
assign MEM[37508] = MEM[17841] + MEM[17851];
assign MEM[37509] = MEM[17844] + MEM[18064];
assign MEM[37510] = MEM[17845] + MEM[17920];
assign MEM[37511] = MEM[17847] + MEM[17867];
assign MEM[37512] = MEM[17853] + MEM[17916];
assign MEM[37513] = MEM[17856] + MEM[17906];
assign MEM[37514] = MEM[17857] + MEM[17881];
assign MEM[37515] = MEM[17858] + MEM[17900];
assign MEM[37516] = MEM[17863] + MEM[17980];
assign MEM[37517] = MEM[17869] + MEM[17879];
assign MEM[37518] = MEM[17870] + MEM[17915];
assign MEM[37519] = MEM[17871] + MEM[17993];
assign MEM[37520] = MEM[17872] + MEM[17887];
assign MEM[37521] = MEM[17876] + MEM[17994];
assign MEM[37522] = MEM[17878] + MEM[17932];
assign MEM[37523] = MEM[17880] + MEM[17965];
assign MEM[37524] = MEM[17883] + MEM[17895];
assign MEM[37525] = MEM[17885] + MEM[18056];
assign MEM[37526] = MEM[17889] + MEM[17908];
assign MEM[37527] = MEM[17891] + MEM[18112];
assign MEM[37528] = MEM[17893] + MEM[17898];
assign MEM[37529] = MEM[17896] + MEM[17917];
assign MEM[37530] = MEM[17897] + MEM[18044];
assign MEM[37531] = MEM[17899] + MEM[18048];
assign MEM[37532] = MEM[17901] + MEM[18012];
assign MEM[37533] = MEM[17904] + MEM[17922];
assign MEM[37534] = MEM[17910] + MEM[17941];
assign MEM[37535] = MEM[17912] + MEM[17956];
assign MEM[37536] = MEM[17914] + MEM[18000];
assign MEM[37537] = MEM[17918] + MEM[17953];
assign MEM[37538] = MEM[17919] + MEM[17964];
assign MEM[37539] = MEM[17924] + MEM[18119];
assign MEM[37540] = MEM[17925] + MEM[17961];
assign MEM[37541] = MEM[17926] + MEM[17929];
assign MEM[37542] = MEM[17927] + MEM[17939];
assign MEM[37543] = MEM[17928] + MEM[17934];
assign MEM[37544] = MEM[17933] + MEM[17947];
assign MEM[37545] = MEM[17936] + MEM[18021];
assign MEM[37546] = MEM[17940] + MEM[18104];
assign MEM[37547] = MEM[17942] + MEM[18163];
assign MEM[37548] = MEM[17943] + MEM[17955];
assign MEM[37549] = MEM[17944] + MEM[17987];
assign MEM[37550] = MEM[17946] + MEM[18002];
assign MEM[37551] = MEM[17949] + MEM[17978];
assign MEM[37552] = MEM[17950] + MEM[17959];
assign MEM[37553] = MEM[17951] + MEM[18029];
assign MEM[37554] = MEM[17952] + MEM[17998];
assign MEM[37555] = MEM[17957] + MEM[17970];
assign MEM[37556] = MEM[17958] + MEM[18072];
assign MEM[37557] = MEM[17962] + MEM[18260];
assign MEM[37558] = MEM[17963] + MEM[17982];
assign MEM[37559] = MEM[17966] + MEM[18003];
assign MEM[37560] = MEM[17967] + MEM[18018];
assign MEM[37561] = MEM[17968] + MEM[18178];
assign MEM[37562] = MEM[17971] + MEM[18006];
assign MEM[37563] = MEM[17972] + MEM[17975];
assign MEM[37564] = MEM[17974] + MEM[18016];
assign MEM[37565] = MEM[17981] + MEM[18181];
assign MEM[37566] = MEM[17983] + MEM[18038];
assign MEM[37567] = MEM[17984] + MEM[18184];
assign MEM[37568] = MEM[17985] + MEM[17990];
assign MEM[37569] = MEM[17986] + MEM[18026];
assign MEM[37570] = MEM[17988] + MEM[18041];
assign MEM[37571] = MEM[17989] + MEM[17995];
assign MEM[37572] = MEM[17999] + MEM[18031];
assign MEM[37573] = MEM[18001] + MEM[18025];
assign MEM[37574] = MEM[18005] + MEM[18014];
assign MEM[37575] = MEM[18008] + MEM[18179];
assign MEM[37576] = MEM[18009] + MEM[18149];
assign MEM[37577] = MEM[18010] + MEM[18213];
assign MEM[37578] = MEM[18011] + MEM[18087];
assign MEM[37579] = MEM[18013] + MEM[18189];
assign MEM[37580] = MEM[18015] + MEM[18039];
assign MEM[37581] = MEM[18019] + MEM[18188];
assign MEM[37582] = MEM[18022] + MEM[18042];
assign MEM[37583] = MEM[18023] + MEM[18098];
assign MEM[37584] = MEM[18024] + MEM[18047];
assign MEM[37585] = MEM[18027] + MEM[18067];
assign MEM[37586] = MEM[18030] + MEM[18106];
assign MEM[37587] = MEM[18032] + MEM[18086];
assign MEM[37588] = MEM[18033] + MEM[18052];
assign MEM[37589] = MEM[18034] + MEM[18201];
assign MEM[37590] = MEM[18035] + MEM[18094];
assign MEM[37591] = MEM[18036] + MEM[18218];
assign MEM[37592] = MEM[18037] + MEM[18125];
assign MEM[37593] = MEM[18040] + MEM[18066];
assign MEM[37594] = MEM[18045] + MEM[18101];
assign MEM[37595] = MEM[18046] + MEM[18153];
assign MEM[37596] = MEM[18050] + MEM[18053];
assign MEM[37597] = MEM[18051] + MEM[18084];
assign MEM[37598] = MEM[18054] + MEM[18071];
assign MEM[37599] = MEM[18055] + MEM[18092];
assign MEM[37600] = MEM[18057] + MEM[18059];
assign MEM[37601] = MEM[18058] + MEM[18141];
assign MEM[37602] = MEM[18060] + MEM[18270];
assign MEM[37603] = MEM[18061] + MEM[18156];
assign MEM[37604] = MEM[18062] + MEM[18111];
assign MEM[37605] = MEM[18063] + MEM[18164];
assign MEM[37606] = MEM[18065] + MEM[18093];
assign MEM[37607] = MEM[18068] + MEM[18571];
assign MEM[37608] = MEM[18070] + MEM[18190];
assign MEM[37609] = MEM[18073] + MEM[18683];
assign MEM[37610] = MEM[18074] + MEM[18161];
assign MEM[37611] = MEM[18075] + MEM[18117];
assign MEM[37612] = MEM[18077] + MEM[18130];
assign MEM[37613] = MEM[18078] + MEM[18083];
assign MEM[37614] = MEM[18080] + MEM[18194];
assign MEM[37615] = MEM[18085] + MEM[18103];
assign MEM[37616] = MEM[18088] + MEM[18176];
assign MEM[37617] = MEM[18090] + MEM[18126];
assign MEM[37618] = MEM[18091] + MEM[18271];
assign MEM[37619] = MEM[18095] + MEM[18105];
assign MEM[37620] = MEM[18096] + MEM[18446];
assign MEM[37621] = MEM[18097] + MEM[18099];
assign MEM[37622] = MEM[18100] + MEM[18136];
assign MEM[37623] = MEM[18107] + MEM[18289];
assign MEM[37624] = MEM[18113] + MEM[18245];
assign MEM[37625] = MEM[18114] + MEM[18131];
assign MEM[37626] = MEM[18115] + MEM[18174];
assign MEM[37627] = MEM[18116] + MEM[18239];
assign MEM[37628] = MEM[18118] + MEM[18152];
assign MEM[37629] = MEM[18121] + MEM[18145];
assign MEM[37630] = MEM[18123] + MEM[18129];
assign MEM[37631] = MEM[18127] + MEM[18187];
assign MEM[37632] = MEM[18128] + MEM[18257];
assign MEM[37633] = MEM[18133] + MEM[18196];
assign MEM[37634] = MEM[18134] + MEM[18250];
assign MEM[37635] = MEM[18135] + MEM[18157];
assign MEM[37636] = MEM[18137] + MEM[18175];
assign MEM[37637] = MEM[18138] + MEM[18282];
assign MEM[37638] = MEM[18140] + MEM[18172];
assign MEM[37639] = MEM[18142] + MEM[18144];
assign MEM[37640] = MEM[18146] + MEM[18202];
assign MEM[37641] = MEM[18150] + MEM[18203];
assign MEM[37642] = MEM[18154] + MEM[18242];
assign MEM[37643] = MEM[18159] + MEM[18323];
assign MEM[37644] = MEM[18160] + MEM[18276];
assign MEM[37645] = MEM[18162] + MEM[18278];
assign MEM[37646] = MEM[18165] + MEM[18227];
assign MEM[37647] = MEM[18167] + MEM[18177];
assign MEM[37648] = MEM[18168] + MEM[18169];
assign MEM[37649] = MEM[18170] + MEM[18273];
assign MEM[37650] = MEM[18171] + MEM[18173];
assign MEM[37651] = MEM[18180] + MEM[18224];
assign MEM[37652] = MEM[18182] + MEM[18186];
assign MEM[37653] = MEM[18185] + MEM[18246];
assign MEM[37654] = MEM[18191] + MEM[18206];
assign MEM[37655] = MEM[18192] + MEM[18216];
assign MEM[37656] = MEM[18193] + MEM[18236];
assign MEM[37657] = MEM[18197] + MEM[18493];
assign MEM[37658] = MEM[18198] + MEM[18208];
assign MEM[37659] = MEM[18199] + MEM[18217];
assign MEM[37660] = MEM[18200] + MEM[18222];
assign MEM[37661] = MEM[18204] + MEM[18251];
assign MEM[37662] = MEM[18205] + MEM[18221];
assign MEM[37663] = MEM[18207] + MEM[18280];
assign MEM[37664] = MEM[18209] + MEM[18212];
assign MEM[37665] = MEM[18211] + MEM[18387];
assign MEM[37666] = MEM[18214] + MEM[18215];
assign MEM[37667] = MEM[18219] + MEM[18269];
assign MEM[37668] = MEM[18220] + MEM[18277];
assign MEM[37669] = MEM[18225] + MEM[18291];
assign MEM[37670] = MEM[18226] + MEM[18349];
assign MEM[37671] = MEM[18228] + MEM[18274];
assign MEM[37672] = MEM[18229] + MEM[18266];
assign MEM[37673] = MEM[18230] + MEM[18304];
assign MEM[37674] = MEM[18232] + MEM[18376];
assign MEM[37675] = MEM[18233] + MEM[18235];
assign MEM[37676] = MEM[18234] + MEM[18341];
assign MEM[37677] = MEM[18237] + MEM[18343];
assign MEM[37678] = MEM[18238] + MEM[18283];
assign MEM[37679] = MEM[18244] + MEM[18346];
assign MEM[37680] = MEM[18247] + MEM[18306];
assign MEM[37681] = MEM[18248] + MEM[18443];
assign MEM[37682] = MEM[18249] + MEM[18478];
assign MEM[37683] = MEM[18252] + MEM[18263];
assign MEM[37684] = MEM[18253] + MEM[18324];
assign MEM[37685] = MEM[18256] + MEM[18264];
assign MEM[37686] = MEM[18259] + MEM[18321];
assign MEM[37687] = MEM[18262] + MEM[18401];
assign MEM[37688] = MEM[18267] + MEM[18362];
assign MEM[37689] = MEM[18268] + MEM[18292];
assign MEM[37690] = MEM[18272] + MEM[18311];
assign MEM[37691] = MEM[18275] + MEM[18285];
assign MEM[37692] = MEM[18279] + MEM[18286];
assign MEM[37693] = MEM[18281] + MEM[18329];
assign MEM[37694] = MEM[18284] + MEM[18293];
assign MEM[37695] = MEM[18287] + MEM[18310];
assign MEM[37696] = MEM[18288] + MEM[18512];
assign MEM[37697] = MEM[18290] + MEM[18412];
assign MEM[37698] = MEM[18294] + MEM[18322];
assign MEM[37699] = MEM[18295] + MEM[18384];
assign MEM[37700] = MEM[18296] + MEM[18348];
assign MEM[37701] = MEM[18297] + MEM[18330];
assign MEM[37702] = MEM[18298] + MEM[18336];
assign MEM[37703] = MEM[18299] + MEM[18339];
assign MEM[37704] = MEM[18300] + MEM[18302];
assign MEM[37705] = MEM[18301] + MEM[18334];
assign MEM[37706] = MEM[18303] + MEM[18386];
assign MEM[37707] = MEM[18305] + MEM[18434];
assign MEM[37708] = MEM[18308] + MEM[18397];
assign MEM[37709] = MEM[18309] + MEM[18375];
assign MEM[37710] = MEM[18312] + MEM[18445];
assign MEM[37711] = MEM[18313] + MEM[18393];
assign MEM[37712] = MEM[18314] + MEM[18415];
assign MEM[37713] = MEM[18317] + MEM[18489];
assign MEM[37714] = MEM[18318] + MEM[18407];
assign MEM[37715] = MEM[18320] + MEM[18369];
assign MEM[37716] = MEM[18326] + MEM[18351];
assign MEM[37717] = MEM[18327] + MEM[18430];
assign MEM[37718] = MEM[18328] + MEM[18360];
assign MEM[37719] = MEM[18331] + MEM[18385];
assign MEM[37720] = MEM[18332] + MEM[18355];
assign MEM[37721] = MEM[18335] + MEM[18418];
assign MEM[37722] = MEM[18337] + MEM[18357];
assign MEM[37723] = MEM[18342] + MEM[18374];
assign MEM[37724] = MEM[18345] + MEM[18356];
assign MEM[37725] = MEM[18347] + MEM[18379];
assign MEM[37726] = MEM[18350] + MEM[18464];
assign MEM[37727] = MEM[18353] + MEM[18382];
assign MEM[37728] = MEM[18354] + MEM[18502];
assign MEM[37729] = MEM[18359] + MEM[18371];
assign MEM[37730] = MEM[18364] + MEM[18435];
assign MEM[37731] = MEM[18365] + MEM[18426];
assign MEM[37732] = MEM[18366] + MEM[18466];
assign MEM[37733] = MEM[18368] + MEM[18377];
assign MEM[37734] = MEM[18370] + MEM[18424];
assign MEM[37735] = MEM[18373] + MEM[18586];
assign MEM[37736] = MEM[18378] + MEM[18530];
assign MEM[37737] = MEM[18380] + MEM[18400];
assign MEM[37738] = MEM[18383] + MEM[18394];
assign MEM[37739] = MEM[18390] + MEM[18440];
assign MEM[37740] = MEM[18392] + MEM[18529];
assign MEM[37741] = MEM[18395] + MEM[18416];
assign MEM[37742] = MEM[18396] + MEM[18458];
assign MEM[37743] = MEM[18398] + MEM[18631];
assign MEM[37744] = MEM[18399] + MEM[18494];
assign MEM[37745] = MEM[18402] + MEM[18422];
assign MEM[37746] = MEM[18403] + MEM[18423];
assign MEM[37747] = MEM[18405] + MEM[18602];
assign MEM[37748] = MEM[18406] + MEM[18451];
assign MEM[37749] = MEM[18409] + MEM[18467];
assign MEM[37750] = MEM[18410] + MEM[18450];
assign MEM[37751] = MEM[18411] + MEM[18477];
assign MEM[37752] = MEM[18414] + MEM[18490];
assign MEM[37753] = MEM[18417] + MEM[18566];
assign MEM[37754] = MEM[18419] + MEM[18439];
assign MEM[37755] = MEM[18420] + MEM[18508];
assign MEM[37756] = MEM[18421] + MEM[18452];
assign MEM[37757] = MEM[18425] + MEM[18455];
assign MEM[37758] = MEM[18427] + MEM[18442];
assign MEM[37759] = MEM[18428] + MEM[18685];
assign MEM[37760] = MEM[18431] + MEM[18531];
assign MEM[37761] = MEM[18432] + MEM[18515];
assign MEM[37762] = MEM[18433] + MEM[18547];
assign MEM[37763] = MEM[18437] + MEM[18660];
assign MEM[37764] = MEM[18448] + MEM[18459];
assign MEM[37765] = MEM[18449] + MEM[18465];
assign MEM[37766] = MEM[18456] + MEM[18575];
assign MEM[37767] = MEM[18460] + MEM[18728];
assign MEM[37768] = MEM[18461] + MEM[18537];
assign MEM[37769] = MEM[18463] + MEM[18501];
assign MEM[37770] = MEM[18468] + MEM[18572];
assign MEM[37771] = MEM[18469] + MEM[18827];
assign MEM[37772] = MEM[18470] + MEM[18475];
assign MEM[37773] = MEM[18471] + MEM[18518];
assign MEM[37774] = MEM[18472] + MEM[18505];
assign MEM[37775] = MEM[18473] + MEM[18497];
assign MEM[37776] = MEM[18479] + MEM[18563];
assign MEM[37777] = MEM[18480] + MEM[18619];
assign MEM[37778] = MEM[18481] + MEM[18533];
assign MEM[37779] = MEM[18482] + MEM[18519];
assign MEM[37780] = MEM[18484] + MEM[18485];
assign MEM[37781] = MEM[18486] + MEM[18487];
assign MEM[37782] = MEM[18488] + MEM[18511];
assign MEM[37783] = MEM[18491] + MEM[18492];
assign MEM[37784] = MEM[18495] + MEM[18513];
assign MEM[37785] = MEM[18496] + MEM[18528];
assign MEM[37786] = MEM[18499] + MEM[18551];
assign MEM[37787] = MEM[18504] + MEM[18627];
assign MEM[37788] = MEM[18506] + MEM[18545];
assign MEM[37789] = MEM[18509] + MEM[18552];
assign MEM[37790] = MEM[18510] + MEM[18764];
assign MEM[37791] = MEM[18514] + MEM[18582];
assign MEM[37792] = MEM[18516] + MEM[18523];
assign MEM[37793] = MEM[18520] + MEM[18535];
assign MEM[37794] = MEM[18522] + MEM[18746];
assign MEM[37795] = MEM[18524] + MEM[18579];
assign MEM[37796] = MEM[18525] + MEM[18532];
assign MEM[37797] = MEM[18527] + MEM[18606];
assign MEM[37798] = MEM[18534] + MEM[18578];
assign MEM[37799] = MEM[18536] + MEM[18541];
assign MEM[37800] = MEM[18538] + MEM[18540];
assign MEM[37801] = MEM[18542] + MEM[18643];
assign MEM[37802] = MEM[18543] + MEM[18562];
assign MEM[37803] = MEM[18544] + MEM[18620];
assign MEM[37804] = MEM[18546] + MEM[18659];
assign MEM[37805] = MEM[18548] + MEM[18597];
assign MEM[37806] = MEM[18549] + MEM[18678];
assign MEM[37807] = MEM[18550] + MEM[18594];
assign MEM[37808] = MEM[18553] + MEM[18748];
assign MEM[37809] = MEM[18555] + MEM[18568];
assign MEM[37810] = MEM[18556] + MEM[18557];
assign MEM[37811] = MEM[18560] + MEM[18603];
assign MEM[37812] = MEM[18561] + MEM[18640];
assign MEM[37813] = MEM[18565] + MEM[18576];
assign MEM[37814] = MEM[18567] + MEM[18625];
assign MEM[37815] = MEM[18570] + MEM[18580];
assign MEM[37816] = MEM[18573] + MEM[18618];
assign MEM[37817] = MEM[18574] + MEM[18706];
assign MEM[37818] = MEM[18577] + MEM[18608];
assign MEM[37819] = MEM[18581] + MEM[18641];
assign MEM[37820] = MEM[18584] + MEM[18585];
assign MEM[37821] = MEM[18587] + MEM[18647];
assign MEM[37822] = MEM[18588] + MEM[18693];
assign MEM[37823] = MEM[18589] + MEM[18677];
assign MEM[37824] = MEM[18592] + MEM[18638];
assign MEM[37825] = MEM[18595] + MEM[18782];
assign MEM[37826] = MEM[18596] + MEM[18730];
assign MEM[37827] = MEM[18600] + MEM[18621];
assign MEM[37828] = MEM[18604] + MEM[18752];
assign MEM[37829] = MEM[18605] + MEM[18615];
assign MEM[37830] = MEM[18611] + MEM[18682];
assign MEM[37831] = MEM[18612] + MEM[18721];
assign MEM[37832] = MEM[18613] + MEM[18668];
assign MEM[37833] = MEM[18614] + MEM[18633];
assign MEM[37834] = MEM[18622] + MEM[18645];
assign MEM[37835] = MEM[18624] + MEM[18727];
assign MEM[37836] = MEM[18626] + MEM[18757];
assign MEM[37837] = MEM[18628] + MEM[18704];
assign MEM[37838] = MEM[18630] + MEM[18713];
assign MEM[37839] = MEM[18632] + MEM[18649];
assign MEM[37840] = MEM[18634] + MEM[18644];
assign MEM[37841] = MEM[18637] + MEM[18665];
assign MEM[37842] = MEM[18639] + MEM[18784];
assign MEM[37843] = MEM[18642] + MEM[18732];
assign MEM[37844] = MEM[18648] + MEM[18662];
assign MEM[37845] = MEM[18650] + MEM[18675];
assign MEM[37846] = MEM[18651] + MEM[18657];
assign MEM[37847] = MEM[18652] + MEM[18821];
assign MEM[37848] = MEM[18653] + MEM[18731];
assign MEM[37849] = MEM[18654] + MEM[18703];
assign MEM[37850] = MEM[18655] + MEM[18658];
assign MEM[37851] = MEM[18656] + MEM[18692];
assign MEM[37852] = MEM[18661] + MEM[18705];
assign MEM[37853] = MEM[18663] + MEM[18822];
assign MEM[37854] = MEM[18666] + MEM[18687];
assign MEM[37855] = MEM[18667] + MEM[18670];
assign MEM[37856] = MEM[18669] + MEM[18707];
assign MEM[37857] = MEM[18671] + MEM[18723];
assign MEM[37858] = MEM[18673] + MEM[18743];
assign MEM[37859] = MEM[18676] + MEM[18733];
assign MEM[37860] = MEM[18679] + MEM[18869];
assign MEM[37861] = MEM[18680] + MEM[18937];
assign MEM[37862] = MEM[18681] + MEM[18871];
assign MEM[37863] = MEM[18684] + MEM[18702];
assign MEM[37864] = MEM[18686] + MEM[18756];
assign MEM[37865] = MEM[18688] + MEM[18774];
assign MEM[37866] = MEM[18690] + MEM[18754];
assign MEM[37867] = MEM[18691] + MEM[18776];
assign MEM[37868] = MEM[18694] + MEM[18722];
assign MEM[37869] = MEM[18695] + MEM[18884];
assign MEM[37870] = MEM[18697] + MEM[18739];
assign MEM[37871] = MEM[18698] + MEM[18744];
assign MEM[37872] = MEM[18699] + MEM[18753];
assign MEM[37873] = MEM[18701] + MEM[18819];
assign MEM[37874] = MEM[18709] + MEM[18726];
assign MEM[37875] = MEM[18710] + MEM[18725];
assign MEM[37876] = MEM[18711] + MEM[18775];
assign MEM[37877] = MEM[18712] + MEM[18887];
assign MEM[37878] = MEM[18714] + MEM[18740];
assign MEM[37879] = MEM[18716] + MEM[18768];
assign MEM[37880] = MEM[18717] + MEM[18829];
assign MEM[37881] = MEM[18719] + MEM[18789];
assign MEM[37882] = MEM[18720] + MEM[18734];
assign MEM[37883] = MEM[18724] + MEM[18826];
assign MEM[37884] = MEM[18729] + MEM[18777];
assign MEM[37885] = MEM[18735] + MEM[18747];
assign MEM[37886] = MEM[18736] + MEM[18769];
assign MEM[37887] = MEM[18737] + MEM[18844];
assign MEM[37888] = MEM[18741] + MEM[18809];
assign MEM[37889] = MEM[18745] + MEM[18876];
assign MEM[37890] = MEM[18749] + MEM[18852];
assign MEM[37891] = MEM[18750] + MEM[19007];
assign MEM[37892] = MEM[18751] + MEM[18766];
assign MEM[37893] = MEM[18755] + MEM[18823];
assign MEM[37894] = MEM[18759] + MEM[18781];
assign MEM[37895] = MEM[18760] + MEM[18934];
assign MEM[37896] = MEM[18761] + MEM[18960];
assign MEM[37897] = MEM[18763] + MEM[18830];
assign MEM[37898] = MEM[18765] + MEM[18818];
assign MEM[37899] = MEM[18767] + MEM[18894];
assign MEM[37900] = MEM[18770] + MEM[18874];
assign MEM[37901] = MEM[18771] + MEM[18801];
assign MEM[37902] = MEM[18778] + MEM[19020];
assign MEM[37903] = MEM[18779] + MEM[18803];
assign MEM[37904] = MEM[18780] + MEM[18802];
assign MEM[37905] = MEM[18783] + MEM[18935];
assign MEM[37906] = MEM[18785] + MEM[18797];
assign MEM[37907] = MEM[18787] + MEM[18998];
assign MEM[37908] = MEM[18788] + MEM[18841];
assign MEM[37909] = MEM[18791] + MEM[18881];
assign MEM[37910] = MEM[18792] + MEM[18904];
assign MEM[37911] = MEM[18793] + MEM[18922];
assign MEM[37912] = MEM[18794] + MEM[18836];
assign MEM[37913] = MEM[18795] + MEM[18843];
assign MEM[37914] = MEM[18796] + MEM[18931];
assign MEM[37915] = MEM[18798] + MEM[18854];
assign MEM[37916] = MEM[18805] + MEM[18817];
assign MEM[37917] = MEM[18806] + MEM[18861];
assign MEM[37918] = MEM[18807] + MEM[18812];
assign MEM[37919] = MEM[18808] + MEM[18865];
assign MEM[37920] = MEM[18811] + MEM[18814];
assign MEM[37921] = MEM[18813] + MEM[18832];
assign MEM[37922] = MEM[18820] + MEM[18842];
assign MEM[37923] = MEM[18828] + MEM[18834];
assign MEM[37924] = MEM[18831] + MEM[18833];
assign MEM[37925] = MEM[18835] + MEM[18864];
assign MEM[37926] = MEM[18837] + MEM[18879];
assign MEM[37927] = MEM[18838] + MEM[18892];
assign MEM[37928] = MEM[18845] + MEM[18853];
assign MEM[37929] = MEM[18847] + MEM[18868];
assign MEM[37930] = MEM[18848] + MEM[18946];
assign MEM[37931] = MEM[18850] + MEM[18867];
assign MEM[37932] = MEM[18851] + MEM[18964];
assign MEM[37933] = MEM[18856] + MEM[18860];
assign MEM[37934] = MEM[18857] + MEM[18872];
assign MEM[37935] = MEM[18858] + MEM[18873];
assign MEM[37936] = MEM[18859] + MEM[18898];
assign MEM[37937] = MEM[18862] + MEM[18878];
assign MEM[37938] = MEM[18866] + MEM[18919];
assign MEM[37939] = MEM[18870] + MEM[18901];
assign MEM[37940] = MEM[18875] + MEM[18897];
assign MEM[37941] = MEM[18877] + MEM[18908];
assign MEM[37942] = MEM[18880] + MEM[18957];
assign MEM[37943] = MEM[18882] + MEM[18890];
assign MEM[37944] = MEM[18883] + MEM[19013];
assign MEM[37945] = MEM[18886] + MEM[18984];
assign MEM[37946] = MEM[18888] + MEM[18914];
assign MEM[37947] = MEM[18889] + MEM[18917];
assign MEM[37948] = MEM[18893] + MEM[18932];
assign MEM[37949] = MEM[18896] + MEM[18930];
assign MEM[37950] = MEM[18900] + MEM[19055];
assign MEM[37951] = MEM[18906] + MEM[18974];
assign MEM[37952] = MEM[18907] + MEM[19133];
assign MEM[37953] = MEM[18909] + MEM[18982];
assign MEM[37954] = MEM[18910] + MEM[18988];
assign MEM[37955] = MEM[18912] + MEM[19064];
assign MEM[37956] = MEM[18913] + MEM[18962];
assign MEM[37957] = MEM[18915] + MEM[18996];
assign MEM[37958] = MEM[18916] + MEM[19002];
assign MEM[37959] = MEM[18918] + MEM[18924];
assign MEM[37960] = MEM[18920] + MEM[18959];
assign MEM[37961] = MEM[18923] + MEM[18981];
assign MEM[37962] = MEM[18925] + MEM[18979];
assign MEM[37963] = MEM[18928] + MEM[18947];
assign MEM[37964] = MEM[18929] + MEM[19158];
assign MEM[37965] = MEM[18933] + MEM[18968];
assign MEM[37966] = MEM[18938] + MEM[18971];
assign MEM[37967] = MEM[18939] + MEM[19088];
assign MEM[37968] = MEM[18940] + MEM[18953];
assign MEM[37969] = MEM[18943] + MEM[18983];
assign MEM[37970] = MEM[18944] + MEM[18965];
assign MEM[37971] = MEM[18945] + MEM[18955];
assign MEM[37972] = MEM[18949] + MEM[19037];
assign MEM[37973] = MEM[18950] + MEM[18992];
assign MEM[37974] = MEM[18951] + MEM[19113];
assign MEM[37975] = MEM[18952] + MEM[19015];
assign MEM[37976] = MEM[18954] + MEM[19009];
assign MEM[37977] = MEM[18961] + MEM[19068];
assign MEM[37978] = MEM[18963] + MEM[19053];
assign MEM[37979] = MEM[18967] + MEM[18980];
assign MEM[37980] = MEM[18969] + MEM[19071];
assign MEM[37981] = MEM[18973] + MEM[19163];
assign MEM[37982] = MEM[18976] + MEM[18989];
assign MEM[37983] = MEM[18977] + MEM[19049];
assign MEM[37984] = MEM[18978] + MEM[19032];
assign MEM[37985] = MEM[18986] + MEM[19067];
assign MEM[37986] = MEM[18990] + MEM[19003];
assign MEM[37987] = MEM[18991] + MEM[19069];
assign MEM[37988] = MEM[18993] + MEM[19026];
assign MEM[37989] = MEM[18994] + MEM[19001];
assign MEM[37990] = MEM[18995] + MEM[19047];
assign MEM[37991] = MEM[18997] + MEM[19264];
assign MEM[37992] = MEM[18999] + MEM[19100];
assign MEM[37993] = MEM[19000] + MEM[19014];
assign MEM[37994] = MEM[19004] + MEM[19056];
assign MEM[37995] = MEM[19006] + MEM[19119];
assign MEM[37996] = MEM[19011] + MEM[19145];
assign MEM[37997] = MEM[19012] + MEM[19094];
assign MEM[37998] = MEM[19016] + MEM[19028];
assign MEM[37999] = MEM[19017] + MEM[19033];
assign MEM[38000] = MEM[19018] + MEM[19063];
assign MEM[38001] = MEM[19019] + MEM[19105];
assign MEM[38002] = MEM[19022] + MEM[19070];
assign MEM[38003] = MEM[19023] + MEM[19058];
assign MEM[38004] = MEM[19024] + MEM[19048];
assign MEM[38005] = MEM[19025] + MEM[19142];
assign MEM[38006] = MEM[19027] + MEM[19135];
assign MEM[38007] = MEM[19029] + MEM[19043];
assign MEM[38008] = MEM[19031] + MEM[19042];
assign MEM[38009] = MEM[19035] + MEM[19107];
assign MEM[38010] = MEM[19036] + MEM[19065];
assign MEM[38011] = MEM[19038] + MEM[19092];
assign MEM[38012] = MEM[19039] + MEM[19080];
assign MEM[38013] = MEM[19041] + MEM[19180];
assign MEM[38014] = MEM[19044] + MEM[19243];
assign MEM[38015] = MEM[19046] + MEM[19141];
assign MEM[38016] = MEM[19050] + MEM[19072];
assign MEM[38017] = MEM[19052] + MEM[19057];
assign MEM[38018] = MEM[19060] + MEM[19115];
assign MEM[38019] = MEM[19062] + MEM[19123];
assign MEM[38020] = MEM[19066] + MEM[19287];
assign MEM[38021] = MEM[19073] + MEM[19118];
assign MEM[38022] = MEM[19074] + MEM[19111];
assign MEM[38023] = MEM[19076] + MEM[19195];
assign MEM[38024] = MEM[19077] + MEM[19184];
assign MEM[38025] = MEM[19078] + MEM[19153];
assign MEM[38026] = MEM[19079] + MEM[19189];
assign MEM[38027] = MEM[19083] + MEM[19097];
assign MEM[38028] = MEM[19084] + MEM[19215];
assign MEM[38029] = MEM[19085] + MEM[19194];
assign MEM[38030] = MEM[19086] + MEM[19387];
assign MEM[38031] = MEM[19087] + MEM[19151];
assign MEM[38032] = MEM[19090] + MEM[19124];
assign MEM[38033] = MEM[19093] + MEM[19245];
assign MEM[38034] = MEM[19095] + MEM[19166];
assign MEM[38035] = MEM[19096] + MEM[19162];
assign MEM[38036] = MEM[19099] + MEM[19103];
assign MEM[38037] = MEM[19101] + MEM[19147];
assign MEM[38038] = MEM[19102] + MEM[19202];
assign MEM[38039] = MEM[19104] + MEM[19137];
assign MEM[38040] = MEM[19106] + MEM[19181];
assign MEM[38041] = MEM[19109] + MEM[19331];
assign MEM[38042] = MEM[19110] + MEM[19301];
assign MEM[38043] = MEM[19112] + MEM[19154];
assign MEM[38044] = MEM[19117] + MEM[19196];
assign MEM[38045] = MEM[19120] + MEM[19122];
assign MEM[38046] = MEM[19121] + MEM[19176];
assign MEM[38047] = MEM[19125] + MEM[19165];
assign MEM[38048] = MEM[19126] + MEM[19168];
assign MEM[38049] = MEM[19127] + MEM[19279];
assign MEM[38050] = MEM[19128] + MEM[19170];
assign MEM[38051] = MEM[19129] + MEM[19132];
assign MEM[38052] = MEM[19131] + MEM[19188];
assign MEM[38053] = MEM[19134] + MEM[19306];
assign MEM[38054] = MEM[19136] + MEM[19167];
assign MEM[38055] = MEM[19138] + MEM[19182];
assign MEM[38056] = MEM[19139] + MEM[19169];
assign MEM[38057] = MEM[19144] + MEM[19173];
assign MEM[38058] = MEM[19146] + MEM[19148];
assign MEM[38059] = MEM[19149] + MEM[19246];
assign MEM[38060] = MEM[19156] + MEM[19157];
assign MEM[38061] = MEM[19159] + MEM[19186];
assign MEM[38062] = MEM[19160] + MEM[19290];
assign MEM[38063] = MEM[19161] + MEM[19259];
assign MEM[38064] = MEM[19164] + MEM[19344];
assign MEM[38065] = MEM[19172] + MEM[19214];
assign MEM[38066] = MEM[19174] + MEM[19523];
assign MEM[38067] = MEM[19175] + MEM[19219];
assign MEM[38068] = MEM[19177] + MEM[19310];
assign MEM[38069] = MEM[19179] + MEM[19221];
assign MEM[38070] = MEM[19185] + MEM[19204];
assign MEM[38071] = MEM[19187] + MEM[19251];
assign MEM[38072] = MEM[19190] + MEM[19234];
assign MEM[38073] = MEM[19191] + MEM[19212];
assign MEM[38074] = MEM[19192] + MEM[19321];
assign MEM[38075] = MEM[19193] + MEM[19520];
assign MEM[38076] = MEM[19197] + MEM[19255];
assign MEM[38077] = MEM[19198] + MEM[19266];
assign MEM[38078] = MEM[19199] + MEM[19289];
assign MEM[38079] = MEM[19200] + MEM[19257];
assign MEM[38080] = MEM[19203] + MEM[19238];
assign MEM[38081] = MEM[19205] + MEM[19299];
assign MEM[38082] = MEM[19206] + MEM[19207];
assign MEM[38083] = MEM[19208] + MEM[19230];
assign MEM[38084] = MEM[19209] + MEM[19253];
assign MEM[38085] = MEM[19210] + MEM[19240];
assign MEM[38086] = MEM[19213] + MEM[19385];
assign MEM[38087] = MEM[19216] + MEM[19293];
assign MEM[38088] = MEM[19217] + MEM[19352];
assign MEM[38089] = MEM[19218] + MEM[19280];
assign MEM[38090] = MEM[19220] + MEM[19313];
assign MEM[38091] = MEM[19222] + MEM[19227];
assign MEM[38092] = MEM[19223] + MEM[19272];
assign MEM[38093] = MEM[19224] + MEM[19231];
assign MEM[38094] = MEM[19229] + MEM[19307];
assign MEM[38095] = MEM[19232] + MEM[19248];
assign MEM[38096] = MEM[19233] + MEM[19496];
assign MEM[38097] = MEM[19235] + MEM[19270];
assign MEM[38098] = MEM[19237] + MEM[19361];
assign MEM[38099] = MEM[19241] + MEM[19332];
assign MEM[38100] = MEM[19249] + MEM[19309];
assign MEM[38101] = MEM[19252] + MEM[19338];
assign MEM[38102] = MEM[19254] + MEM[19452];
assign MEM[38103] = MEM[19256] + MEM[19334];
assign MEM[38104] = MEM[19258] + MEM[19378];
assign MEM[38105] = MEM[19261] + MEM[19380];
assign MEM[38106] = MEM[19262] + MEM[19267];
assign MEM[38107] = MEM[19265] + MEM[19354];
assign MEM[38108] = MEM[19268] + MEM[19295];
assign MEM[38109] = MEM[19269] + MEM[19285];
assign MEM[38110] = MEM[19273] + MEM[19277];
assign MEM[38111] = MEM[19274] + MEM[19291];
assign MEM[38112] = MEM[19278] + MEM[19416];
assign MEM[38113] = MEM[19281] + MEM[19316];
assign MEM[38114] = MEM[19282] + MEM[19345];
assign MEM[38115] = MEM[19284] + MEM[19360];
assign MEM[38116] = MEM[19286] + MEM[19297];
assign MEM[38117] = MEM[19288] + MEM[19324];
assign MEM[38118] = MEM[19292] + MEM[19405];
assign MEM[38119] = MEM[19294] + MEM[19322];
assign MEM[38120] = MEM[19298] + MEM[19339];
assign MEM[38121] = MEM[19300] + MEM[19311];
assign MEM[38122] = MEM[19302] + MEM[19394];
assign MEM[38123] = MEM[19303] + MEM[19349];
assign MEM[38124] = MEM[19304] + MEM[19379];
assign MEM[38125] = MEM[19305] + MEM[19358];
assign MEM[38126] = MEM[19308] + MEM[19340];
assign MEM[38127] = MEM[19312] + MEM[19367];
assign MEM[38128] = MEM[19314] + MEM[19315];
assign MEM[38129] = MEM[19317] + MEM[19366];
assign MEM[38130] = MEM[19318] + MEM[19368];
assign MEM[38131] = MEM[19323] + MEM[19363];
assign MEM[38132] = MEM[19325] + MEM[19330];
assign MEM[38133] = MEM[19326] + MEM[19327];
assign MEM[38134] = MEM[19328] + MEM[19364];
assign MEM[38135] = MEM[19329] + MEM[19577];
assign MEM[38136] = MEM[19333] + MEM[19373];
assign MEM[38137] = MEM[19335] + MEM[19443];
assign MEM[38138] = MEM[19337] + MEM[19469];
assign MEM[38139] = MEM[19346] + MEM[19390];
assign MEM[38140] = MEM[19347] + MEM[19362];
assign MEM[38141] = MEM[19348] + MEM[19474];
assign MEM[38142] = MEM[19350] + MEM[19433];
assign MEM[38143] = MEM[19351] + MEM[19388];
assign MEM[38144] = MEM[19353] + MEM[19459];
assign MEM[38145] = MEM[19356] + MEM[19365];
assign MEM[38146] = MEM[19369] + MEM[19485];
assign MEM[38147] = MEM[19370] + MEM[19386];
assign MEM[38148] = MEM[19372] + MEM[19615];
assign MEM[38149] = MEM[19374] + MEM[19454];
assign MEM[38150] = MEM[19375] + MEM[19381];
assign MEM[38151] = MEM[19376] + MEM[19626];
assign MEM[38152] = MEM[19377] + MEM[19424];
assign MEM[38153] = MEM[19383] + MEM[19438];
assign MEM[38154] = MEM[19384] + MEM[19428];
assign MEM[38155] = MEM[19389] + MEM[19398];
assign MEM[38156] = MEM[19391] + MEM[19447];
assign MEM[38157] = MEM[19392] + MEM[19508];
assign MEM[38158] = MEM[19393] + MEM[19440];
assign MEM[38159] = MEM[19396] + MEM[19429];
assign MEM[38160] = MEM[19397] + MEM[19449];
assign MEM[38161] = MEM[19399] + MEM[19402];
assign MEM[38162] = MEM[19400] + MEM[19413];
assign MEM[38163] = MEM[19401] + MEM[19467];
assign MEM[38164] = MEM[19404] + MEM[19490];
assign MEM[38165] = MEM[19406] + MEM[19605];
assign MEM[38166] = MEM[19407] + MEM[19503];
assign MEM[38167] = MEM[19408] + MEM[19484];
assign MEM[38168] = MEM[19410] + MEM[19458];
assign MEM[38169] = MEM[19411] + MEM[19422];
assign MEM[38170] = MEM[19417] + MEM[19494];
assign MEM[38171] = MEM[19418] + MEM[19426];
assign MEM[38172] = MEM[19419] + MEM[19617];
assign MEM[38173] = MEM[19420] + MEM[19547];
assign MEM[38174] = MEM[19421] + MEM[19480];
assign MEM[38175] = MEM[19423] + MEM[19560];
assign MEM[38176] = MEM[19427] + MEM[19608];
assign MEM[38177] = MEM[19430] + MEM[19552];
assign MEM[38178] = MEM[19432] + MEM[19435];
assign MEM[38179] = MEM[19434] + MEM[19534];
assign MEM[38180] = MEM[19436] + MEM[19791];
assign MEM[38181] = MEM[19442] + MEM[19509];
assign MEM[38182] = MEM[19444] + MEM[19512];
assign MEM[38183] = MEM[19446] + MEM[19519];
assign MEM[38184] = MEM[19448] + MEM[19549];
assign MEM[38185] = MEM[19450] + MEM[19527];
assign MEM[38186] = MEM[19451] + MEM[19461];
assign MEM[38187] = MEM[19453] + MEM[19460];
assign MEM[38188] = MEM[19455] + MEM[19457];
assign MEM[38189] = MEM[19456] + MEM[19696];
assign MEM[38190] = MEM[19462] + MEM[19650];
assign MEM[38191] = MEM[19464] + MEM[19539];
assign MEM[38192] = MEM[19465] + MEM[19504];
assign MEM[38193] = MEM[19466] + MEM[19489];
assign MEM[38194] = MEM[19468] + MEM[19510];
assign MEM[38195] = MEM[19470] + MEM[19473];
assign MEM[38196] = MEM[19471] + MEM[19528];
assign MEM[38197] = MEM[19472] + MEM[19488];
assign MEM[38198] = MEM[19475] + MEM[19515];
assign MEM[38199] = MEM[19476] + MEM[19517];
assign MEM[38200] = MEM[19477] + MEM[19533];
assign MEM[38201] = MEM[19481] + MEM[19498];
assign MEM[38202] = MEM[19486] + MEM[19499];
assign MEM[38203] = MEM[19491] + MEM[19501];
assign MEM[38204] = MEM[19492] + MEM[19537];
assign MEM[38205] = MEM[19493] + MEM[19532];
assign MEM[38206] = MEM[19495] + MEM[19595];
assign MEM[38207] = MEM[19500] + MEM[19548];
assign MEM[38208] = MEM[19502] + MEM[19563];
assign MEM[38209] = MEM[19505] + MEM[19614];
assign MEM[38210] = MEM[19506] + MEM[19590];
assign MEM[38211] = MEM[19507] + MEM[19550];
assign MEM[38212] = MEM[19511] + MEM[19542];
assign MEM[38213] = MEM[19513] + MEM[19538];
assign MEM[38214] = MEM[19514] + MEM[19647];
assign MEM[38215] = MEM[19516] + MEM[19568];
assign MEM[38216] = MEM[19518] + MEM[19584];
assign MEM[38217] = MEM[19521] + MEM[19708];
assign MEM[38218] = MEM[19522] + MEM[19663];
assign MEM[38219] = MEM[19524] + MEM[19661];
assign MEM[38220] = MEM[19525] + MEM[19541];
assign MEM[38221] = MEM[19526] + MEM[19624];
assign MEM[38222] = MEM[19529] + MEM[19720];
assign MEM[38223] = MEM[19530] + MEM[19635];
assign MEM[38224] = MEM[19531] + MEM[19633];
assign MEM[38225] = MEM[19536] + MEM[19555];
assign MEM[38226] = MEM[19540] + MEM[19606];
assign MEM[38227] = MEM[19543] + MEM[19616];
assign MEM[38228] = MEM[19544] + MEM[19567];
assign MEM[38229] = MEM[19546] + MEM[19593];
assign MEM[38230] = MEM[19551] + MEM[19620];
assign MEM[38231] = MEM[19553] + MEM[19586];
assign MEM[38232] = MEM[19556] + MEM[19582];
assign MEM[38233] = MEM[19557] + MEM[19632];
assign MEM[38234] = MEM[19559] + MEM[19666];
assign MEM[38235] = MEM[19561] + MEM[20107];
assign MEM[38236] = MEM[19562] + MEM[19613];
assign MEM[38237] = MEM[19565] + MEM[19703];
assign MEM[38238] = MEM[19569] + MEM[19594];
assign MEM[38239] = MEM[19570] + MEM[19648];
assign MEM[38240] = MEM[19571] + MEM[19643];
assign MEM[38241] = MEM[19572] + MEM[19746];
assign MEM[38242] = MEM[19574] + MEM[19714];
assign MEM[38243] = MEM[19576] + MEM[19676];
assign MEM[38244] = MEM[19578] + MEM[19580];
assign MEM[38245] = MEM[19581] + MEM[19641];
assign MEM[38246] = MEM[19583] + MEM[19602];
assign MEM[38247] = MEM[19587] + MEM[19655];
assign MEM[38248] = MEM[19589] + MEM[19630];
assign MEM[38249] = MEM[19591] + MEM[19660];
assign MEM[38250] = MEM[19592] + MEM[19680];
assign MEM[38251] = MEM[19597] + MEM[19598];
assign MEM[38252] = MEM[19599] + MEM[19609];
assign MEM[38253] = MEM[19601] + MEM[19611];
assign MEM[38254] = MEM[19603] + MEM[19625];
assign MEM[38255] = MEM[19607] + MEM[19687];
assign MEM[38256] = MEM[19610] + MEM[19712];
assign MEM[38257] = MEM[19612] + MEM[19767];
assign MEM[38258] = MEM[19618] + MEM[19744];
assign MEM[38259] = MEM[19619] + MEM[19622];
assign MEM[38260] = MEM[19621] + MEM[19652];
assign MEM[38261] = MEM[19627] + MEM[19631];
assign MEM[38262] = MEM[19629] + MEM[19684];
assign MEM[38263] = MEM[19634] + MEM[19734];
assign MEM[38264] = MEM[19636] + MEM[19669];
assign MEM[38265] = MEM[19640] + MEM[19654];
assign MEM[38266] = MEM[19644] + MEM[19873];
assign MEM[38267] = MEM[19646] + MEM[19697];
assign MEM[38268] = MEM[19649] + MEM[19694];
assign MEM[38269] = MEM[19651] + MEM[19754];
assign MEM[38270] = MEM[19653] + MEM[19670];
assign MEM[38271] = MEM[19657] + MEM[19686];
assign MEM[38272] = MEM[19658] + MEM[19682];
assign MEM[38273] = MEM[19662] + MEM[19679];
assign MEM[38274] = MEM[19664] + MEM[19711];
assign MEM[38275] = MEM[19665] + MEM[19769];
assign MEM[38276] = MEM[19667] + MEM[19727];
assign MEM[38277] = MEM[19668] + MEM[19776];
assign MEM[38278] = MEM[19671] + MEM[19883];
assign MEM[38279] = MEM[19673] + MEM[19713];
assign MEM[38280] = MEM[19674] + MEM[19729];
assign MEM[38281] = MEM[19675] + MEM[19692];
assign MEM[38282] = MEM[19678] + MEM[19707];
assign MEM[38283] = MEM[19681] + MEM[19704];
assign MEM[38284] = MEM[19683] + MEM[19733];
assign MEM[38285] = MEM[19685] + MEM[19737];
assign MEM[38286] = MEM[19688] + MEM[19775];
assign MEM[38287] = MEM[19691] + MEM[19840];
assign MEM[38288] = MEM[19695] + MEM[19702];
assign MEM[38289] = MEM[19698] + MEM[19830];
assign MEM[38290] = MEM[19699] + MEM[19805];
assign MEM[38291] = MEM[19701] + MEM[19725];
assign MEM[38292] = MEM[19709] + MEM[19722];
assign MEM[38293] = MEM[19710] + MEM[19850];
assign MEM[38294] = MEM[19715] + MEM[19750];
assign MEM[38295] = MEM[19716] + MEM[19788];
assign MEM[38296] = MEM[19717] + MEM[19766];
assign MEM[38297] = MEM[19718] + MEM[19763];
assign MEM[38298] = MEM[19719] + MEM[19726];
assign MEM[38299] = MEM[19721] + MEM[19863];
assign MEM[38300] = MEM[19723] + MEM[19825];
assign MEM[38301] = MEM[19728] + MEM[19741];
assign MEM[38302] = MEM[19730] + MEM[19901];
assign MEM[38303] = MEM[19731] + MEM[19836];
assign MEM[38304] = MEM[19732] + MEM[19795];
assign MEM[38305] = MEM[19735] + MEM[19761];
assign MEM[38306] = MEM[19736] + MEM[19748];
assign MEM[38307] = MEM[19738] + MEM[19773];
assign MEM[38308] = MEM[19740] + MEM[19777];
assign MEM[38309] = MEM[19742] + MEM[20106];
assign MEM[38310] = MEM[19745] + MEM[19839];
assign MEM[38311] = MEM[19747] + MEM[19841];
assign MEM[38312] = MEM[19749] + MEM[19782];
assign MEM[38313] = MEM[19751] + MEM[19760];
assign MEM[38314] = MEM[19752] + MEM[19857];
assign MEM[38315] = MEM[19753] + MEM[19755];
assign MEM[38316] = MEM[19756] + MEM[19774];
assign MEM[38317] = MEM[19757] + MEM[19933];
assign MEM[38318] = MEM[19758] + MEM[19855];
assign MEM[38319] = MEM[19759] + MEM[19871];
assign MEM[38320] = MEM[19762] + MEM[19851];
assign MEM[38321] = MEM[19765] + MEM[19804];
assign MEM[38322] = MEM[19768] + MEM[19824];
assign MEM[38323] = MEM[19770] + MEM[19780];
assign MEM[38324] = MEM[19771] + MEM[19816];
assign MEM[38325] = MEM[19772] + MEM[19809];
assign MEM[38326] = MEM[19778] + MEM[19779];
assign MEM[38327] = MEM[19781] + MEM[19807];
assign MEM[38328] = MEM[19783] + MEM[19962];
assign MEM[38329] = MEM[19784] + MEM[19800];
assign MEM[38330] = MEM[19785] + MEM[19786];
assign MEM[38331] = MEM[19790] + MEM[19808];
assign MEM[38332] = MEM[19792] + MEM[19903];
assign MEM[38333] = MEM[19793] + MEM[19812];
assign MEM[38334] = MEM[19794] + MEM[19953];
assign MEM[38335] = MEM[19797] + MEM[19942];
assign MEM[38336] = MEM[19798] + MEM[19818];
assign MEM[38337] = MEM[19802] + MEM[19912];
assign MEM[38338] = MEM[19810] + MEM[19862];
assign MEM[38339] = MEM[19813] + MEM[19980];
assign MEM[38340] = MEM[19814] + MEM[19864];
assign MEM[38341] = MEM[19815] + MEM[19834];
assign MEM[38342] = MEM[19817] + MEM[19899];
assign MEM[38343] = MEM[19819] + MEM[19833];
assign MEM[38344] = MEM[19820] + MEM[19996];
assign MEM[38345] = MEM[19822] + MEM[19860];
assign MEM[38346] = MEM[19826] + MEM[19898];
assign MEM[38347] = MEM[19827] + MEM[19894];
assign MEM[38348] = MEM[19829] + MEM[19881];
assign MEM[38349] = MEM[19831] + MEM[20077];
assign MEM[38350] = MEM[19842] + MEM[19943];
assign MEM[38351] = MEM[19844] + MEM[19906];
assign MEM[38352] = MEM[19845] + MEM[19847];
assign MEM[38353] = MEM[19849] + MEM[19985];
assign MEM[38354] = MEM[19852] + MEM[19891];
assign MEM[38355] = MEM[19853] + MEM[19885];
assign MEM[38356] = MEM[19854] + MEM[19911];
assign MEM[38357] = MEM[19858] + MEM[19893];
assign MEM[38358] = MEM[19859] + MEM[19966];
assign MEM[38359] = MEM[19861] + MEM[19877];
assign MEM[38360] = MEM[19866] + MEM[19867];
assign MEM[38361] = MEM[19868] + MEM[20117];
assign MEM[38362] = MEM[19869] + MEM[20010];
assign MEM[38363] = MEM[19870] + MEM[19905];
assign MEM[38364] = MEM[19872] + MEM[19874];
assign MEM[38365] = MEM[19875] + MEM[19890];
assign MEM[38366] = MEM[19876] + MEM[19910];
assign MEM[38367] = MEM[19879] + MEM[19917];
assign MEM[38368] = MEM[19882] + MEM[20019];
assign MEM[38369] = MEM[19884] + MEM[19989];
assign MEM[38370] = MEM[19887] + MEM[19960];
assign MEM[38371] = MEM[19888] + MEM[19947];
assign MEM[38372] = MEM[19889] + MEM[19957];
assign MEM[38373] = MEM[19892] + MEM[19934];
assign MEM[38374] = MEM[19896] + MEM[19925];
assign MEM[38375] = MEM[19897] + MEM[19930];
assign MEM[38376] = MEM[19904] + MEM[20025];
assign MEM[38377] = MEM[19907] + MEM[19954];
assign MEM[38378] = MEM[19908] + MEM[19939];
assign MEM[38379] = MEM[19909] + MEM[19941];
assign MEM[38380] = MEM[19913] + MEM[19927];
assign MEM[38381] = MEM[19914] + MEM[19987];
assign MEM[38382] = MEM[19918] + MEM[19970];
assign MEM[38383] = MEM[19919] + MEM[19983];
assign MEM[38384] = MEM[19920] + MEM[20054];
assign MEM[38385] = MEM[19921] + MEM[19971];
assign MEM[38386] = MEM[19922] + MEM[19997];
assign MEM[38387] = MEM[19923] + MEM[19952];
assign MEM[38388] = MEM[19924] + MEM[20072];
assign MEM[38389] = MEM[19928] + MEM[19959];
assign MEM[38390] = MEM[19929] + MEM[20091];
assign MEM[38391] = MEM[19931] + MEM[19955];
assign MEM[38392] = MEM[19932] + MEM[20070];
assign MEM[38393] = MEM[19935] + MEM[20095];
assign MEM[38394] = MEM[19936] + MEM[19945];
assign MEM[38395] = MEM[19937] + MEM[19979];
assign MEM[38396] = MEM[19938] + MEM[19946];
assign MEM[38397] = MEM[19940] + MEM[20006];
assign MEM[38398] = MEM[19944] + MEM[20055];
assign MEM[38399] = MEM[19949] + MEM[20002];
assign MEM[38400] = MEM[19951] + MEM[19964];
assign MEM[38401] = MEM[19958] + MEM[19978];
assign MEM[38402] = MEM[19963] + MEM[20125];
assign MEM[38403] = MEM[19965] + MEM[20038];
assign MEM[38404] = MEM[19967] + MEM[19969];
assign MEM[38405] = MEM[19968] + MEM[20012];
assign MEM[38406] = MEM[19973] + MEM[20027];
assign MEM[38407] = MEM[19974] + MEM[20143];
assign MEM[38408] = MEM[19975] + MEM[20016];
assign MEM[38409] = MEM[19976] + MEM[20008];
assign MEM[38410] = MEM[19977] + MEM[19990];
assign MEM[38411] = MEM[19981] + MEM[20103];
assign MEM[38412] = MEM[19982] + MEM[20051];
assign MEM[38413] = MEM[19986] + MEM[20000];
assign MEM[38414] = MEM[19988] + MEM[19993];
assign MEM[38415] = MEM[19991] + MEM[20206];
assign MEM[38416] = MEM[19992] + MEM[20067];
assign MEM[38417] = MEM[19995] + MEM[20022];
assign MEM[38418] = MEM[19999] + MEM[20013];
assign MEM[38419] = MEM[20001] + MEM[20015];
assign MEM[38420] = MEM[20003] + MEM[20062];
assign MEM[38421] = MEM[20004] + MEM[20042];
assign MEM[38422] = MEM[20005] + MEM[20044];
assign MEM[38423] = MEM[20007] + MEM[20142];
assign MEM[38424] = MEM[20009] + MEM[20087];
assign MEM[38425] = MEM[20011] + MEM[20024];
assign MEM[38426] = MEM[20014] + MEM[20083];
assign MEM[38427] = MEM[20018] + MEM[20030];
assign MEM[38428] = MEM[20020] + MEM[20086];
assign MEM[38429] = MEM[20023] + MEM[20115];
assign MEM[38430] = MEM[20026] + MEM[20047];
assign MEM[38431] = MEM[20028] + MEM[20177];
assign MEM[38432] = MEM[20031] + MEM[20060];
assign MEM[38433] = MEM[20032] + MEM[20040];
assign MEM[38434] = MEM[20034] + MEM[20075];
assign MEM[38435] = MEM[20036] + MEM[20049];
assign MEM[38436] = MEM[20037] + MEM[20123];
assign MEM[38437] = MEM[20039] + MEM[20116];
assign MEM[38438] = MEM[20041] + MEM[20045];
assign MEM[38439] = MEM[20043] + MEM[20113];
assign MEM[38440] = MEM[20048] + MEM[20241];
assign MEM[38441] = MEM[20050] + MEM[20098];
assign MEM[38442] = MEM[20052] + MEM[20074];
assign MEM[38443] = MEM[20053] + MEM[20079];
assign MEM[38444] = MEM[20058] + MEM[20063];
assign MEM[38445] = MEM[20064] + MEM[20144];
assign MEM[38446] = MEM[20065] + MEM[20089];
assign MEM[38447] = MEM[20068] + MEM[20088];
assign MEM[38448] = MEM[20071] + MEM[20112];
assign MEM[38449] = MEM[20073] + MEM[20084];
assign MEM[38450] = MEM[20076] + MEM[20226];
assign MEM[38451] = MEM[20078] + MEM[20141];
assign MEM[38452] = MEM[20080] + MEM[20104];
assign MEM[38453] = MEM[20081] + MEM[20255];
assign MEM[38454] = MEM[20082] + MEM[20111];
assign MEM[38455] = MEM[20092] + MEM[20152];
assign MEM[38456] = MEM[20093] + MEM[20097];
assign MEM[38457] = MEM[20094] + MEM[20119];
assign MEM[38458] = MEM[20096] + MEM[20151];
assign MEM[38459] = MEM[20099] + MEM[20158];
assign MEM[38460] = MEM[20100] + MEM[20170];
assign MEM[38461] = MEM[20101] + MEM[20155];
assign MEM[38462] = MEM[20102] + MEM[20129];
assign MEM[38463] = MEM[20105] + MEM[20162];
assign MEM[38464] = MEM[20108] + MEM[20227];
assign MEM[38465] = MEM[20109] + MEM[20295];
assign MEM[38466] = MEM[20110] + MEM[20261];
assign MEM[38467] = MEM[20114] + MEM[20120];
assign MEM[38468] = MEM[20121] + MEM[20252];
assign MEM[38469] = MEM[20124] + MEM[20173];
assign MEM[38470] = MEM[20126] + MEM[20482];
assign MEM[38471] = MEM[20127] + MEM[20332];
assign MEM[38472] = MEM[20128] + MEM[20197];
assign MEM[38473] = MEM[20132] + MEM[20273];
assign MEM[38474] = MEM[20133] + MEM[20192];
assign MEM[38475] = MEM[20134] + MEM[20337];
assign MEM[38476] = MEM[20135] + MEM[20230];
assign MEM[38477] = MEM[20136] + MEM[20307];
assign MEM[38478] = MEM[20137] + MEM[20163];
assign MEM[38479] = MEM[20138] + MEM[20237];
assign MEM[38480] = MEM[20139] + MEM[20275];
assign MEM[38481] = MEM[20140] + MEM[20156];
assign MEM[38482] = MEM[20145] + MEM[20214];
assign MEM[38483] = MEM[20146] + MEM[20529];
assign MEM[38484] = MEM[20148] + MEM[20205];
assign MEM[38485] = MEM[20149] + MEM[20293];
assign MEM[38486] = MEM[20153] + MEM[20234];
assign MEM[38487] = MEM[20154] + MEM[20180];
assign MEM[38488] = MEM[20157] + MEM[20165];
assign MEM[38489] = MEM[20159] + MEM[20213];
assign MEM[38490] = MEM[20160] + MEM[20408];
assign MEM[38491] = MEM[20161] + MEM[20185];
assign MEM[38492] = MEM[20164] + MEM[20184];
assign MEM[38493] = MEM[20166] + MEM[20181];
assign MEM[38494] = MEM[20167] + MEM[20208];
assign MEM[38495] = MEM[20169] + MEM[20178];
assign MEM[38496] = MEM[20171] + MEM[20179];
assign MEM[38497] = MEM[20172] + MEM[20201];
assign MEM[38498] = MEM[20174] + MEM[20232];
assign MEM[38499] = MEM[20175] + MEM[20196];
assign MEM[38500] = MEM[20182] + MEM[20291];
assign MEM[38501] = MEM[20183] + MEM[20198];
assign MEM[38502] = MEM[20187] + MEM[20415];
assign MEM[38503] = MEM[20188] + MEM[20248];
assign MEM[38504] = MEM[20190] + MEM[20203];
assign MEM[38505] = MEM[20191] + MEM[20264];
assign MEM[38506] = MEM[20193] + MEM[20253];
assign MEM[38507] = MEM[20194] + MEM[20279];
assign MEM[38508] = MEM[20195] + MEM[20256];
assign MEM[38509] = MEM[20199] + MEM[20454];
assign MEM[38510] = MEM[20200] + MEM[20409];
assign MEM[38511] = MEM[20207] + MEM[20346];
assign MEM[38512] = MEM[20209] + MEM[20328];
assign MEM[38513] = MEM[20210] + MEM[20285];
assign MEM[38514] = MEM[20211] + MEM[20453];
assign MEM[38515] = MEM[20212] + MEM[20235];
assign MEM[38516] = MEM[20216] + MEM[20238];
assign MEM[38517] = MEM[20217] + MEM[20243];
assign MEM[38518] = MEM[20219] + MEM[20246];
assign MEM[38519] = MEM[20220] + MEM[20229];
assign MEM[38520] = MEM[20223] + MEM[20371];
assign MEM[38521] = MEM[20224] + MEM[20348];
assign MEM[38522] = MEM[20228] + MEM[20263];
assign MEM[38523] = MEM[20231] + MEM[20254];
assign MEM[38524] = MEM[20233] + MEM[20289];
assign MEM[38525] = MEM[20239] + MEM[20520];
assign MEM[38526] = MEM[20249] + MEM[20276];
assign MEM[38527] = MEM[20250] + MEM[20303];
assign MEM[38528] = MEM[20251] + MEM[20298];
assign MEM[38529] = MEM[20257] + MEM[20266];
assign MEM[38530] = MEM[20258] + MEM[20320];
assign MEM[38531] = MEM[20260] + MEM[20323];
assign MEM[38532] = MEM[20262] + MEM[20286];
assign MEM[38533] = MEM[20267] + MEM[20403];
assign MEM[38534] = MEM[20268] + MEM[20302];
assign MEM[38535] = MEM[20269] + MEM[20548];
assign MEM[38536] = MEM[20270] + MEM[20305];
assign MEM[38537] = MEM[20272] + MEM[20308];
assign MEM[38538] = MEM[20277] + MEM[20324];
assign MEM[38539] = MEM[20281] + MEM[20315];
assign MEM[38540] = MEM[20282] + MEM[20327];
assign MEM[38541] = MEM[20283] + MEM[20427];
assign MEM[38542] = MEM[20284] + MEM[20416];
assign MEM[38543] = MEM[20287] + MEM[20354];
assign MEM[38544] = MEM[20288] + MEM[20361];
assign MEM[38545] = MEM[20290] + MEM[20301];
assign MEM[38546] = MEM[20292] + MEM[20383];
assign MEM[38547] = MEM[20296] + MEM[20336];
assign MEM[38548] = MEM[20299] + MEM[20310];
assign MEM[38549] = MEM[20300] + MEM[20333];
assign MEM[38550] = MEM[20306] + MEM[20313];
assign MEM[38551] = MEM[20309] + MEM[20343];
assign MEM[38552] = MEM[20311] + MEM[20352];
assign MEM[38553] = MEM[20312] + MEM[20340];
assign MEM[38554] = MEM[20316] + MEM[20425];
assign MEM[38555] = MEM[20317] + MEM[20339];
assign MEM[38556] = MEM[20318] + MEM[20469];
assign MEM[38557] = MEM[20319] + MEM[20331];
assign MEM[38558] = MEM[20321] + MEM[20329];
assign MEM[38559] = MEM[20322] + MEM[20670];
assign MEM[38560] = MEM[20326] + MEM[20461];
assign MEM[38561] = MEM[20330] + MEM[20367];
assign MEM[38562] = MEM[20334] + MEM[20477];
assign MEM[38563] = MEM[20335] + MEM[20412];
assign MEM[38564] = MEM[20338] + MEM[20370];
assign MEM[38565] = MEM[20341] + MEM[20496];
assign MEM[38566] = MEM[20342] + MEM[20381];
assign MEM[38567] = MEM[20344] + MEM[20420];
assign MEM[38568] = MEM[20347] + MEM[20385];
assign MEM[38569] = MEM[20350] + MEM[20391];
assign MEM[38570] = MEM[20353] + MEM[20504];
assign MEM[38571] = MEM[20356] + MEM[20511];
assign MEM[38572] = MEM[20357] + MEM[20399];
assign MEM[38573] = MEM[20358] + MEM[20365];
assign MEM[38574] = MEM[20359] + MEM[20426];
assign MEM[38575] = MEM[20360] + MEM[20404];
assign MEM[38576] = MEM[20362] + MEM[20380];
assign MEM[38577] = MEM[20364] + MEM[20700];
assign MEM[38578] = MEM[20366] + MEM[20500];
assign MEM[38579] = MEM[20368] + MEM[20444];
assign MEM[38580] = MEM[20369] + MEM[20379];
assign MEM[38581] = MEM[20374] + MEM[20392];
assign MEM[38582] = MEM[20375] + MEM[20448];
assign MEM[38583] = MEM[20377] + MEM[20423];
assign MEM[38584] = MEM[20378] + MEM[20601];
assign MEM[38585] = MEM[20382] + MEM[20582];
assign MEM[38586] = MEM[20384] + MEM[20396];
assign MEM[38587] = MEM[20386] + MEM[20443];
assign MEM[38588] = MEM[20387] + MEM[20397];
assign MEM[38589] = MEM[20388] + MEM[20476];
assign MEM[38590] = MEM[20389] + MEM[20432];
assign MEM[38591] = MEM[20390] + MEM[20720];
assign MEM[38592] = MEM[20393] + MEM[20506];
assign MEM[38593] = MEM[20394] + MEM[20411];
assign MEM[38594] = MEM[20395] + MEM[20451];
assign MEM[38595] = MEM[20398] + MEM[20431];
assign MEM[38596] = MEM[20400] + MEM[20472];
assign MEM[38597] = MEM[20401] + MEM[20555];
assign MEM[38598] = MEM[20402] + MEM[20471];
assign MEM[38599] = MEM[20405] + MEM[20459];
assign MEM[38600] = MEM[20406] + MEM[20458];
assign MEM[38601] = MEM[20407] + MEM[20502];
assign MEM[38602] = MEM[20410] + MEM[20583];
assign MEM[38603] = MEM[20413] + MEM[20577];
assign MEM[38604] = MEM[20417] + MEM[20537];
assign MEM[38605] = MEM[20418] + MEM[20445];
assign MEM[38606] = MEM[20419] + MEM[20532];
assign MEM[38607] = MEM[20424] + MEM[20648];
assign MEM[38608] = MEM[20429] + MEM[20534];
assign MEM[38609] = MEM[20430] + MEM[20437];
assign MEM[38610] = MEM[20434] + MEM[20447];
assign MEM[38611] = MEM[20435] + MEM[20450];
assign MEM[38612] = MEM[20436] + MEM[20510];
assign MEM[38613] = MEM[20438] + MEM[20462];
assign MEM[38614] = MEM[20439] + MEM[20449];
assign MEM[38615] = MEM[20440] + MEM[20475];
assign MEM[38616] = MEM[20442] + MEM[20483];
assign MEM[38617] = MEM[20452] + MEM[20468];
assign MEM[38618] = MEM[20456] + MEM[20517];
assign MEM[38619] = MEM[20463] + MEM[20589];
assign MEM[38620] = MEM[20464] + MEM[20597];
assign MEM[38621] = MEM[20465] + MEM[20588];
assign MEM[38622] = MEM[20466] + MEM[20569];
assign MEM[38623] = MEM[20467] + MEM[20522];
assign MEM[38624] = MEM[20470] + MEM[20474];
assign MEM[38625] = MEM[20479] + MEM[20632];
assign MEM[38626] = MEM[20484] + MEM[20515];
assign MEM[38627] = MEM[20485] + MEM[20591];
assign MEM[38628] = MEM[20486] + MEM[20599];
assign MEM[38629] = MEM[20487] + MEM[20505];
assign MEM[38630] = MEM[20488] + MEM[20530];
assign MEM[38631] = MEM[20489] + MEM[20493];
assign MEM[38632] = MEM[20490] + MEM[20531];
assign MEM[38633] = MEM[20492] + MEM[20499];
assign MEM[38634] = MEM[20497] + MEM[20628];
assign MEM[38635] = MEM[20498] + MEM[20525];
assign MEM[38636] = MEM[20501] + MEM[20646];
assign MEM[38637] = MEM[20503] + MEM[20549];
assign MEM[38638] = MEM[20507] + MEM[20523];
assign MEM[38639] = MEM[20509] + MEM[20633];
assign MEM[38640] = MEM[20512] + MEM[20556];
assign MEM[38641] = MEM[20513] + MEM[20624];
assign MEM[38642] = MEM[20514] + MEM[20613];
assign MEM[38643] = MEM[20518] + MEM[20746];
assign MEM[38644] = MEM[20519] + MEM[20546];
assign MEM[38645] = MEM[20524] + MEM[20621];
assign MEM[38646] = MEM[20526] + MEM[20551];
assign MEM[38647] = MEM[20527] + MEM[20607];
assign MEM[38648] = MEM[20528] + MEM[20554];
assign MEM[38649] = MEM[20533] + MEM[20641];
assign MEM[38650] = MEM[20538] + MEM[20587];
assign MEM[38651] = MEM[20539] + MEM[20545];
assign MEM[38652] = MEM[20540] + MEM[20600];
assign MEM[38653] = MEM[20541] + MEM[20604];
assign MEM[38654] = MEM[20542] + MEM[20580];
assign MEM[38655] = MEM[20543] + MEM[20818];
assign MEM[38656] = MEM[20544] + MEM[20943];
assign MEM[38657] = MEM[20552] + MEM[20667];
assign MEM[38658] = MEM[20553] + MEM[20572];
assign MEM[38659] = MEM[20560] + MEM[20570];
assign MEM[38660] = MEM[20562] + MEM[20719];
assign MEM[38661] = MEM[20563] + MEM[20565];
assign MEM[38662] = MEM[20564] + MEM[20658];
assign MEM[38663] = MEM[20566] + MEM[20611];
assign MEM[38664] = MEM[20567] + MEM[20702];
assign MEM[38665] = MEM[20568] + MEM[20573];
assign MEM[38666] = MEM[20571] + MEM[20687];
assign MEM[38667] = MEM[20574] + MEM[20704];
assign MEM[38668] = MEM[20576] + MEM[20740];
assign MEM[38669] = MEM[20578] + MEM[20627];
assign MEM[38670] = MEM[20579] + MEM[20837];
assign MEM[38671] = MEM[20581] + MEM[20586];
assign MEM[38672] = MEM[20585] + MEM[20661];
assign MEM[38673] = MEM[20590] + MEM[20631];
assign MEM[38674] = MEM[20593] + MEM[20623];
assign MEM[38675] = MEM[20594] + MEM[20757];
assign MEM[38676] = MEM[20595] + MEM[20731];
assign MEM[38677] = MEM[20596] + MEM[20643];
assign MEM[38678] = MEM[20602] + MEM[20614];
assign MEM[38679] = MEM[20603] + MEM[20722];
assign MEM[38680] = MEM[20605] + MEM[20659];
assign MEM[38681] = MEM[20606] + MEM[20651];
assign MEM[38682] = MEM[20608] + MEM[20642];
assign MEM[38683] = MEM[20610] + MEM[20615];
assign MEM[38684] = MEM[20612] + MEM[20710];
assign MEM[38685] = MEM[20616] + MEM[20685];
assign MEM[38686] = MEM[20617] + MEM[20650];
assign MEM[38687] = MEM[20618] + MEM[20805];
assign MEM[38688] = MEM[20619] + MEM[20666];
assign MEM[38689] = MEM[20620] + MEM[20675];
assign MEM[38690] = MEM[20625] + MEM[20779];
assign MEM[38691] = MEM[20626] + MEM[20688];
assign MEM[38692] = MEM[20629] + MEM[20679];
assign MEM[38693] = MEM[20630] + MEM[20663];
assign MEM[38694] = MEM[20634] + MEM[20712];
assign MEM[38695] = MEM[20635] + MEM[20878];
assign MEM[38696] = MEM[20636] + MEM[20981];
assign MEM[38697] = MEM[20637] + MEM[20652];
assign MEM[38698] = MEM[20638] + MEM[20645];
assign MEM[38699] = MEM[20639] + MEM[20707];
assign MEM[38700] = MEM[20644] + MEM[20751];
assign MEM[38701] = MEM[20647] + MEM[20715];
assign MEM[38702] = MEM[20653] + MEM[20787];
assign MEM[38703] = MEM[20654] + MEM[20655];
assign MEM[38704] = MEM[20656] + MEM[20717];
assign MEM[38705] = MEM[20660] + MEM[20781];
assign MEM[38706] = MEM[20662] + MEM[20674];
assign MEM[38707] = MEM[20665] + MEM[20684];
assign MEM[38708] = MEM[20668] + MEM[20997];
assign MEM[38709] = MEM[20669] + MEM[20806];
assign MEM[38710] = MEM[20672] + MEM[20725];
assign MEM[38711] = MEM[20676] + MEM[20690];
assign MEM[38712] = MEM[20677] + MEM[20750];
assign MEM[38713] = MEM[20678] + MEM[20758];
assign MEM[38714] = MEM[20680] + MEM[20769];
assign MEM[38715] = MEM[20683] + MEM[20718];
assign MEM[38716] = MEM[20686] + MEM[20695];
assign MEM[38717] = MEM[20689] + MEM[20705];
assign MEM[38718] = MEM[20691] + MEM[20789];
assign MEM[38719] = MEM[20692] + MEM[20728];
assign MEM[38720] = MEM[20698] + MEM[20738];
assign MEM[38721] = MEM[20708] + MEM[20713];
assign MEM[38722] = MEM[20709] + MEM[20721];
assign MEM[38723] = MEM[20711] + MEM[20867];
assign MEM[38724] = MEM[20723] + MEM[20734];
assign MEM[38725] = MEM[20724] + MEM[20832];
assign MEM[38726] = MEM[20726] + MEM[20822];
assign MEM[38727] = MEM[20727] + MEM[20791];
assign MEM[38728] = MEM[20729] + MEM[20875];
assign MEM[38729] = MEM[20730] + MEM[20760];
assign MEM[38730] = MEM[20732] + MEM[20748];
assign MEM[38731] = MEM[20733] + MEM[21028];
assign MEM[38732] = MEM[20735] + MEM[20754];
assign MEM[38733] = MEM[20736] + MEM[20767];
assign MEM[38734] = MEM[20739] + MEM[20942];
assign MEM[38735] = MEM[20741] + MEM[20743];
assign MEM[38736] = MEM[20744] + MEM[20788];
assign MEM[38737] = MEM[20745] + MEM[20829];
assign MEM[38738] = MEM[20747] + MEM[20824];
assign MEM[38739] = MEM[20753] + MEM[20759];
assign MEM[38740] = MEM[20755] + MEM[20964];
assign MEM[38741] = MEM[20756] + MEM[20859];
assign MEM[38742] = MEM[20762] + MEM[20800];
assign MEM[38743] = MEM[20763] + MEM[20796];
assign MEM[38744] = MEM[20766] + MEM[20783];
assign MEM[38745] = MEM[20771] + MEM[20905];
assign MEM[38746] = MEM[20773] + MEM[20949];
assign MEM[38747] = MEM[20774] + MEM[20790];
assign MEM[38748] = MEM[20776] + MEM[20853];
assign MEM[38749] = MEM[20777] + MEM[20846];
assign MEM[38750] = MEM[20778] + MEM[20793];
assign MEM[38751] = MEM[20792] + MEM[20920];
assign MEM[38752] = MEM[20794] + MEM[20866];
assign MEM[38753] = MEM[20797] + MEM[20918];
assign MEM[38754] = MEM[20798] + MEM[20885];
assign MEM[38755] = MEM[20799] + MEM[21189];
assign MEM[38756] = MEM[20801] + MEM[20892];
assign MEM[38757] = MEM[20802] + MEM[20830];
assign MEM[38758] = MEM[20803] + MEM[21312];
assign MEM[38759] = MEM[20804] + MEM[20820];
assign MEM[38760] = MEM[20807] + MEM[20907];
assign MEM[38761] = MEM[20808] + MEM[20958];
assign MEM[38762] = MEM[20809] + MEM[20882];
assign MEM[38763] = MEM[20810] + MEM[20915];
assign MEM[38764] = MEM[20811] + MEM[20821];
assign MEM[38765] = MEM[20813] + MEM[20836];
assign MEM[38766] = MEM[20814] + MEM[20926];
assign MEM[38767] = MEM[20816] + MEM[20917];
assign MEM[38768] = MEM[20819] + MEM[20826];
assign MEM[38769] = MEM[20823] + MEM[20844];
assign MEM[38770] = MEM[20825] + MEM[21254];
assign MEM[38771] = MEM[20827] + MEM[20833];
assign MEM[38772] = MEM[20828] + MEM[20843];
assign MEM[38773] = MEM[20834] + MEM[20894];
assign MEM[38774] = MEM[20835] + MEM[20887];
assign MEM[38775] = MEM[20838] + MEM[20855];
assign MEM[38776] = MEM[20839] + MEM[20888];
assign MEM[38777] = MEM[20840] + MEM[20856];
assign MEM[38778] = MEM[20841] + MEM[20881];
assign MEM[38779] = MEM[20842] + MEM[20899];
assign MEM[38780] = MEM[20848] + MEM[20903];
assign MEM[38781] = MEM[20849] + MEM[20941];
assign MEM[38782] = MEM[20850] + MEM[21176];
assign MEM[38783] = MEM[20851] + MEM[20950];
assign MEM[38784] = MEM[20852] + MEM[21129];
assign MEM[38785] = MEM[20854] + MEM[20862];
assign MEM[38786] = MEM[20861] + MEM[20924];
assign MEM[38787] = MEM[20864] + MEM[21144];
assign MEM[38788] = MEM[20865] + MEM[21001];
assign MEM[38789] = MEM[20868] + MEM[20896];
assign MEM[38790] = MEM[20869] + MEM[20939];
assign MEM[38791] = MEM[20870] + MEM[20976];
assign MEM[38792] = MEM[20871] + MEM[20901];
assign MEM[38793] = MEM[20872] + MEM[20884];
assign MEM[38794] = MEM[20873] + MEM[20910];
assign MEM[38795] = MEM[20874] + MEM[20931];
assign MEM[38796] = MEM[20876] + MEM[20945];
assign MEM[38797] = MEM[20877] + MEM[20879];
assign MEM[38798] = MEM[20883] + MEM[20963];
assign MEM[38799] = MEM[20886] + MEM[20889];
assign MEM[38800] = MEM[20891] + MEM[21018];
assign MEM[38801] = MEM[20895] + MEM[20948];
assign MEM[38802] = MEM[20897] + MEM[20912];
assign MEM[38803] = MEM[20898] + MEM[20902];
assign MEM[38804] = MEM[20900] + MEM[20904];
assign MEM[38805] = MEM[20906] + MEM[20967];
assign MEM[38806] = MEM[20908] + MEM[20980];
assign MEM[38807] = MEM[20909] + MEM[20928];
assign MEM[38808] = MEM[20911] + MEM[20987];
assign MEM[38809] = MEM[20913] + MEM[20922];
assign MEM[38810] = MEM[20914] + MEM[20940];
assign MEM[38811] = MEM[20919] + MEM[21048];
assign MEM[38812] = MEM[20925] + MEM[21262];
assign MEM[38813] = MEM[20927] + MEM[20947];
assign MEM[38814] = MEM[20929] + MEM[20937];
assign MEM[38815] = MEM[20930] + MEM[20960];
assign MEM[38816] = MEM[20932] + MEM[20953];
assign MEM[38817] = MEM[20934] + MEM[20973];
assign MEM[38818] = MEM[20935] + MEM[21000];
assign MEM[38819] = MEM[20936] + MEM[20996];
assign MEM[38820] = MEM[20938] + MEM[20977];
assign MEM[38821] = MEM[20944] + MEM[21077];
assign MEM[38822] = MEM[20946] + MEM[21038];
assign MEM[38823] = MEM[20951] + MEM[20966];
assign MEM[38824] = MEM[20952] + MEM[20959];
assign MEM[38825] = MEM[20956] + MEM[21047];
assign MEM[38826] = MEM[20957] + MEM[21030];
assign MEM[38827] = MEM[20961] + MEM[20999];
assign MEM[38828] = MEM[20962] + MEM[21014];
assign MEM[38829] = MEM[20968] + MEM[21019];
assign MEM[38830] = MEM[20969] + MEM[20985];
assign MEM[38831] = MEM[20970] + MEM[21169];
assign MEM[38832] = MEM[20971] + MEM[21302];
assign MEM[38833] = MEM[20972] + MEM[21031];
assign MEM[38834] = MEM[20975] + MEM[21002];
assign MEM[38835] = MEM[20978] + MEM[21175];
assign MEM[38836] = MEM[20979] + MEM[21194];
assign MEM[38837] = MEM[20982] + MEM[21004];
assign MEM[38838] = MEM[20983] + MEM[21051];
assign MEM[38839] = MEM[20984] + MEM[21105];
assign MEM[38840] = MEM[20986] + MEM[21011];
assign MEM[38841] = MEM[20988] + MEM[21010];
assign MEM[38842] = MEM[20989] + MEM[20992];
assign MEM[38843] = MEM[20990] + MEM[20991];
assign MEM[38844] = MEM[20993] + MEM[21089];
assign MEM[38845] = MEM[20994] + MEM[21163];
assign MEM[38846] = MEM[20995] + MEM[21053];
assign MEM[38847] = MEM[20998] + MEM[21072];
assign MEM[38848] = MEM[21003] + MEM[21071];
assign MEM[38849] = MEM[21005] + MEM[21020];
assign MEM[38850] = MEM[21006] + MEM[21062];
assign MEM[38851] = MEM[21008] + MEM[21017];
assign MEM[38852] = MEM[21009] + MEM[21021];
assign MEM[38853] = MEM[21012] + MEM[21118];
assign MEM[38854] = MEM[21013] + MEM[21083];
assign MEM[38855] = MEM[21015] + MEM[21114];
assign MEM[38856] = MEM[21016] + MEM[21130];
assign MEM[38857] = MEM[21022] + MEM[21064];
assign MEM[38858] = MEM[21023] + MEM[21251];
assign MEM[38859] = MEM[21024] + MEM[21088];
assign MEM[38860] = MEM[21025] + MEM[21085];
assign MEM[38861] = MEM[21029] + MEM[21140];
assign MEM[38862] = MEM[21032] + MEM[21068];
assign MEM[38863] = MEM[21033] + MEM[21065];
assign MEM[38864] = MEM[21034] + MEM[21125];
assign MEM[38865] = MEM[21035] + MEM[21036];
assign MEM[38866] = MEM[21039] + MEM[21041];
assign MEM[38867] = MEM[21040] + MEM[21073];
assign MEM[38868] = MEM[21042] + MEM[21337];
assign MEM[38869] = MEM[21043] + MEM[21097];
assign MEM[38870] = MEM[21044] + MEM[21075];
assign MEM[38871] = MEM[21045] + MEM[21121];
assign MEM[38872] = MEM[21046] + MEM[21049];
assign MEM[38873] = MEM[21050] + MEM[21134];
assign MEM[38874] = MEM[21052] + MEM[21326];
assign MEM[38875] = MEM[21054] + MEM[21087];
assign MEM[38876] = MEM[21056] + MEM[21106];
assign MEM[38877] = MEM[21057] + MEM[21112];
assign MEM[38878] = MEM[21059] + MEM[21128];
assign MEM[38879] = MEM[21060] + MEM[21093];
assign MEM[38880] = MEM[21063] + MEM[21137];
assign MEM[38881] = MEM[21069] + MEM[21132];
assign MEM[38882] = MEM[21074] + MEM[21243];
assign MEM[38883] = MEM[21078] + MEM[21162];
assign MEM[38884] = MEM[21079] + MEM[21099];
assign MEM[38885] = MEM[21080] + MEM[21359];
assign MEM[38886] = MEM[21081] + MEM[21235];
assign MEM[38887] = MEM[21084] + MEM[21086];
assign MEM[38888] = MEM[21090] + MEM[21101];
assign MEM[38889] = MEM[21092] + MEM[21135];
assign MEM[38890] = MEM[21094] + MEM[21113];
assign MEM[38891] = MEM[21098] + MEM[21119];
assign MEM[38892] = MEM[21102] + MEM[21178];
assign MEM[38893] = MEM[21109] + MEM[21197];
assign MEM[38894] = MEM[21111] + MEM[21196];
assign MEM[38895] = MEM[21115] + MEM[21157];
assign MEM[38896] = MEM[21116] + MEM[21203];
assign MEM[38897] = MEM[21117] + MEM[21138];
assign MEM[38898] = MEM[21120] + MEM[21139];
assign MEM[38899] = MEM[21122] + MEM[21124];
assign MEM[38900] = MEM[21123] + MEM[21160];
assign MEM[38901] = MEM[21126] + MEM[21240];
assign MEM[38902] = MEM[21131] + MEM[21231];
assign MEM[38903] = MEM[21133] + MEM[21154];
assign MEM[38904] = MEM[21141] + MEM[21241];
assign MEM[38905] = MEM[21142] + MEM[21269];
assign MEM[38906] = MEM[21143] + MEM[21388];
assign MEM[38907] = MEM[21145] + MEM[21267];
assign MEM[38908] = MEM[21146] + MEM[21258];
assign MEM[38909] = MEM[21147] + MEM[21182];
assign MEM[38910] = MEM[21148] + MEM[21150];
assign MEM[38911] = MEM[21149] + MEM[21206];
assign MEM[38912] = MEM[21151] + MEM[21156];
assign MEM[38913] = MEM[21152] + MEM[21174];
assign MEM[38914] = MEM[21153] + MEM[21223];
assign MEM[38915] = MEM[21155] + MEM[21172];
assign MEM[38916] = MEM[21158] + MEM[21187];
assign MEM[38917] = MEM[21159] + MEM[21161];
assign MEM[38918] = MEM[21165] + MEM[21301];
assign MEM[38919] = MEM[21166] + MEM[21344];
assign MEM[38920] = MEM[21167] + MEM[21215];
assign MEM[38921] = MEM[21168] + MEM[21479];
assign MEM[38922] = MEM[21170] + MEM[21211];
assign MEM[38923] = MEM[21171] + MEM[21362];
assign MEM[38924] = MEM[21173] + MEM[21191];
assign MEM[38925] = MEM[21177] + MEM[21201];
assign MEM[38926] = MEM[21179] + MEM[21213];
assign MEM[38927] = MEM[21180] + MEM[21199];
assign MEM[38928] = MEM[21183] + MEM[21268];
assign MEM[38929] = MEM[21184] + MEM[21316];
assign MEM[38930] = MEM[21186] + MEM[21271];
assign MEM[38931] = MEM[21188] + MEM[21314];
assign MEM[38932] = MEM[21190] + MEM[21288];
assign MEM[38933] = MEM[21192] + MEM[21214];
assign MEM[38934] = MEM[21193] + MEM[21207];
assign MEM[38935] = MEM[21198] + MEM[21321];
assign MEM[38936] = MEM[21200] + MEM[21205];
assign MEM[38937] = MEM[21202] + MEM[21366];
assign MEM[38938] = MEM[21204] + MEM[21272];
assign MEM[38939] = MEM[21208] + MEM[21274];
assign MEM[38940] = MEM[21209] + MEM[21368];
assign MEM[38941] = MEM[21216] + MEM[21405];
assign MEM[38942] = MEM[21217] + MEM[21393];
assign MEM[38943] = MEM[21218] + MEM[21292];
assign MEM[38944] = MEM[21220] + MEM[21239];
assign MEM[38945] = MEM[21221] + MEM[21352];
assign MEM[38946] = MEM[21222] + MEM[21249];
assign MEM[38947] = MEM[21224] + MEM[21233];
assign MEM[38948] = MEM[21225] + MEM[21336];
assign MEM[38949] = MEM[21226] + MEM[21232];
assign MEM[38950] = MEM[21228] + MEM[21230];
assign MEM[38951] = MEM[21234] + MEM[21285];
assign MEM[38952] = MEM[21237] + MEM[21273];
assign MEM[38953] = MEM[21238] + MEM[21377];
assign MEM[38954] = MEM[21244] + MEM[21252];
assign MEM[38955] = MEM[21245] + MEM[21310];
assign MEM[38956] = MEM[21246] + MEM[21277];
assign MEM[38957] = MEM[21247] + MEM[21281];
assign MEM[38958] = MEM[21250] + MEM[21290];
assign MEM[38959] = MEM[21253] + MEM[21474];
assign MEM[38960] = MEM[21256] + MEM[21309];
assign MEM[38961] = MEM[21257] + MEM[21367];
assign MEM[38962] = MEM[21259] + MEM[21327];
assign MEM[38963] = MEM[21261] + MEM[21275];
assign MEM[38964] = MEM[21263] + MEM[21476];
assign MEM[38965] = MEM[21265] + MEM[21413];
assign MEM[38966] = MEM[21266] + MEM[21497];
assign MEM[38967] = MEM[21270] + MEM[21382];
assign MEM[38968] = MEM[21276] + MEM[21284];
assign MEM[38969] = MEM[21278] + MEM[21451];
assign MEM[38970] = MEM[21279] + MEM[21298];
assign MEM[38971] = MEM[21280] + MEM[21297];
assign MEM[38972] = MEM[21282] + MEM[21318];
assign MEM[38973] = MEM[21283] + MEM[21399];
assign MEM[38974] = MEM[21286] + MEM[21328];
assign MEM[38975] = MEM[21287] + MEM[21320];
assign MEM[38976] = MEM[21289] + MEM[21385];
assign MEM[38977] = MEM[21291] + MEM[21358];
assign MEM[38978] = MEM[21293] + MEM[21317];
assign MEM[38979] = MEM[21299] + MEM[21345];
assign MEM[38980] = MEM[21300] + MEM[21374];
assign MEM[38981] = MEM[21306] + MEM[21414];
assign MEM[38982] = MEM[21308] + MEM[21403];
assign MEM[38983] = MEM[21315] + MEM[21391];
assign MEM[38984] = MEM[21319] + MEM[21499];
assign MEM[38985] = MEM[21323] + MEM[21355];
assign MEM[38986] = MEM[21325] + MEM[21349];
assign MEM[38987] = MEM[21330] + MEM[21389];
assign MEM[38988] = MEM[21332] + MEM[21375];
assign MEM[38989] = MEM[21333] + MEM[21378];
assign MEM[38990] = MEM[21334] + MEM[21365];
assign MEM[38991] = MEM[21335] + MEM[21369];
assign MEM[38992] = MEM[21338] + MEM[21347];
assign MEM[38993] = MEM[21339] + MEM[21492];
assign MEM[38994] = MEM[21340] + MEM[21357];
assign MEM[38995] = MEM[21342] + MEM[21452];
assign MEM[38996] = MEM[21343] + MEM[21503];
assign MEM[38997] = MEM[21346] + MEM[21409];
assign MEM[38998] = MEM[21350] + MEM[21379];
assign MEM[38999] = MEM[21351] + MEM[21356];
assign MEM[39000] = MEM[21360] + MEM[21401];
assign MEM[39001] = MEM[21361] + MEM[21395];
assign MEM[39002] = MEM[21364] + MEM[21614];
assign MEM[39003] = MEM[21370] + MEM[21415];
assign MEM[39004] = MEM[21373] + MEM[21472];
assign MEM[39005] = MEM[21380] + MEM[21563];
assign MEM[39006] = MEM[21383] + MEM[21423];
assign MEM[39007] = MEM[21384] + MEM[21398];
assign MEM[39008] = MEM[21387] + MEM[21443];
assign MEM[39009] = MEM[21390] + MEM[21481];
assign MEM[39010] = MEM[21392] + MEM[21461];
assign MEM[39011] = MEM[21396] + MEM[21468];
assign MEM[39012] = MEM[21397] + MEM[21438];
assign MEM[39013] = MEM[21400] + MEM[21432];
assign MEM[39014] = MEM[21402] + MEM[21450];
assign MEM[39015] = MEM[21406] + MEM[21425];
assign MEM[39016] = MEM[21407] + MEM[21477];
assign MEM[39017] = MEM[21408] + MEM[21434];
assign MEM[39018] = MEM[21410] + MEM[21487];
assign MEM[39019] = MEM[21411] + MEM[21433];
assign MEM[39020] = MEM[21412] + MEM[21490];
assign MEM[39021] = MEM[21416] + MEM[21541];
assign MEM[39022] = MEM[21417] + MEM[21548];
assign MEM[39023] = MEM[21419] + MEM[21576];
assign MEM[39024] = MEM[21420] + MEM[21448];
assign MEM[39025] = MEM[21421] + MEM[21464];
assign MEM[39026] = MEM[21422] + MEM[21446];
assign MEM[39027] = MEM[21424] + MEM[21549];
assign MEM[39028] = MEM[21426] + MEM[21524];
assign MEM[39029] = MEM[21427] + MEM[21471];
assign MEM[39030] = MEM[21429] + MEM[21431];
assign MEM[39031] = MEM[21435] + MEM[21442];
assign MEM[39032] = MEM[21437] + MEM[21639];
assign MEM[39033] = MEM[21439] + MEM[21545];
assign MEM[39034] = MEM[21440] + MEM[21666];
assign MEM[39035] = MEM[21441] + MEM[21648];
assign MEM[39036] = MEM[21444] + MEM[21661];
assign MEM[39037] = MEM[21447] + MEM[21501];
assign MEM[39038] = MEM[21454] + MEM[21515];
assign MEM[39039] = MEM[21455] + MEM[21456];
assign MEM[39040] = MEM[21458] + MEM[21508];
assign MEM[39041] = MEM[21459] + MEM[21725];
assign MEM[39042] = MEM[21460] + MEM[21525];
assign MEM[39043] = MEM[21462] + MEM[21523];
assign MEM[39044] = MEM[21466] + MEM[21467];
assign MEM[39045] = MEM[21469] + MEM[21506];
assign MEM[39046] = MEM[21470] + MEM[21537];
assign MEM[39047] = MEM[21475] + MEM[21603];
assign MEM[39048] = MEM[21478] + MEM[21533];
assign MEM[39049] = MEM[21480] + MEM[21496];
assign MEM[39050] = MEM[21482] + MEM[21527];
assign MEM[39051] = MEM[21483] + MEM[21539];
assign MEM[39052] = MEM[21485] + MEM[21671];
assign MEM[39053] = MEM[21486] + MEM[21489];
assign MEM[39054] = MEM[21488] + MEM[21587];
assign MEM[39055] = MEM[21491] + MEM[21498];
assign MEM[39056] = MEM[21493] + MEM[21553];
assign MEM[39057] = MEM[21494] + MEM[21572];
assign MEM[39058] = MEM[21495] + MEM[21677];
assign MEM[39059] = MEM[21500] + MEM[21514];
assign MEM[39060] = MEM[21502] + MEM[21560];
assign MEM[39061] = MEM[21505] + MEM[21636];
assign MEM[39062] = MEM[21507] + MEM[21577];
assign MEM[39063] = MEM[21509] + MEM[21518];
assign MEM[39064] = MEM[21511] + MEM[21829];
assign MEM[39065] = MEM[21512] + MEM[21551];
assign MEM[39066] = MEM[21513] + MEM[21662];
assign MEM[39067] = MEM[21516] + MEM[21651];
assign MEM[39068] = MEM[21519] + MEM[21668];
assign MEM[39069] = MEM[21520] + MEM[21542];
assign MEM[39070] = MEM[21521] + MEM[21609];
assign MEM[39071] = MEM[21522] + MEM[21540];
assign MEM[39072] = MEM[21526] + MEM[21566];
assign MEM[39073] = MEM[21528] + MEM[21637];
assign MEM[39074] = MEM[21529] + MEM[21716];
assign MEM[39075] = MEM[21531] + MEM[21728];
assign MEM[39076] = MEM[21532] + MEM[21626];
assign MEM[39077] = MEM[21534] + MEM[21634];
assign MEM[39078] = MEM[21535] + MEM[21559];
assign MEM[39079] = MEM[21543] + MEM[21564];
assign MEM[39080] = MEM[21544] + MEM[21569];
assign MEM[39081] = MEM[21546] + MEM[21891];
assign MEM[39082] = MEM[21550] + MEM[21555];
assign MEM[39083] = MEM[21552] + MEM[21594];
assign MEM[39084] = MEM[21554] + MEM[21621];
assign MEM[39085] = MEM[21556] + MEM[21573];
assign MEM[39086] = MEM[21557] + MEM[21608];
assign MEM[39087] = MEM[21561] + MEM[21664];
assign MEM[39088] = MEM[21562] + MEM[21610];
assign MEM[39089] = MEM[21565] + MEM[21601];
assign MEM[39090] = MEM[21567] + MEM[21653];
assign MEM[39091] = MEM[21568] + MEM[21586];
assign MEM[39092] = MEM[21574] + MEM[21616];
assign MEM[39093] = MEM[21575] + MEM[21593];
assign MEM[39094] = MEM[21578] + MEM[21679];
assign MEM[39095] = MEM[21579] + MEM[21743];
assign MEM[39096] = MEM[21580] + MEM[21591];
assign MEM[39097] = MEM[21582] + MEM[21655];
assign MEM[39098] = MEM[21583] + MEM[21602];
assign MEM[39099] = MEM[21584] + MEM[21612];
assign MEM[39100] = MEM[21585] + MEM[21665];
assign MEM[39101] = MEM[21588] + MEM[21729];
assign MEM[39102] = MEM[21589] + MEM[21599];
assign MEM[39103] = MEM[21592] + MEM[21604];
assign MEM[39104] = MEM[21597] + MEM[21710];
assign MEM[39105] = MEM[21600] + MEM[21684];
assign MEM[39106] = MEM[21605] + MEM[21795];
assign MEM[39107] = MEM[21606] + MEM[21617];
assign MEM[39108] = MEM[21611] + MEM[21660];
assign MEM[39109] = MEM[21613] + MEM[21846];
assign MEM[39110] = MEM[21615] + MEM[21654];
assign MEM[39111] = MEM[21619] + MEM[21656];
assign MEM[39112] = MEM[21620] + MEM[21705];
assign MEM[39113] = MEM[21622] + MEM[21742];
assign MEM[39114] = MEM[21623] + MEM[21817];
assign MEM[39115] = MEM[21624] + MEM[21779];
assign MEM[39116] = MEM[21625] + MEM[21789];
assign MEM[39117] = MEM[21628] + MEM[21658];
assign MEM[39118] = MEM[21629] + MEM[21764];
assign MEM[39119] = MEM[21630] + MEM[21635];
assign MEM[39120] = MEM[21631] + MEM[21745];
assign MEM[39121] = MEM[21632] + MEM[21703];
assign MEM[39122] = MEM[21638] + MEM[21650];
assign MEM[39123] = MEM[21641] + MEM[21682];
assign MEM[39124] = MEM[21643] + MEM[21657];
assign MEM[39125] = MEM[21644] + MEM[21678];
assign MEM[39126] = MEM[21646] + MEM[21681];
assign MEM[39127] = MEM[21649] + MEM[21794];
assign MEM[39128] = MEM[21652] + MEM[21726];
assign MEM[39129] = MEM[21659] + MEM[21688];
assign MEM[39130] = MEM[21663] + MEM[21747];
assign MEM[39131] = MEM[21667] + MEM[21757];
assign MEM[39132] = MEM[21669] + MEM[21778];
assign MEM[39133] = MEM[21670] + MEM[22032];
assign MEM[39134] = MEM[21672] + MEM[21706];
assign MEM[39135] = MEM[21673] + MEM[21699];
assign MEM[39136] = MEM[21674] + MEM[21719];
assign MEM[39137] = MEM[21675] + MEM[21689];
assign MEM[39138] = MEM[21676] + MEM[21723];
assign MEM[39139] = MEM[21680] + MEM[21709];
assign MEM[39140] = MEM[21685] + MEM[21690];
assign MEM[39141] = MEM[21686] + MEM[21746];
assign MEM[39142] = MEM[21691] + MEM[21980];
assign MEM[39143] = MEM[21692] + MEM[21926];
assign MEM[39144] = MEM[21693] + MEM[21768];
assign MEM[39145] = MEM[21694] + MEM[21696];
assign MEM[39146] = MEM[21695] + MEM[21875];
assign MEM[39147] = MEM[21697] + MEM[21708];
assign MEM[39148] = MEM[21698] + MEM[21751];
assign MEM[39149] = MEM[21700] + MEM[21786];
assign MEM[39150] = MEM[21701] + MEM[21803];
assign MEM[39151] = MEM[21702] + MEM[21758];
assign MEM[39152] = MEM[21704] + MEM[21836];
assign MEM[39153] = MEM[21707] + MEM[21711];
assign MEM[39154] = MEM[21712] + MEM[21812];
assign MEM[39155] = MEM[21714] + MEM[21735];
assign MEM[39156] = MEM[21715] + MEM[21763];
assign MEM[39157] = MEM[21717] + MEM[21910];
assign MEM[39158] = MEM[21720] + MEM[21734];
assign MEM[39159] = MEM[21721] + MEM[21756];
assign MEM[39160] = MEM[21727] + MEM[21759];
assign MEM[39161] = MEM[21730] + MEM[21854];
assign MEM[39162] = MEM[21733] + MEM[21775];
assign MEM[39163] = MEM[21736] + MEM[21807];
assign MEM[39164] = MEM[21737] + MEM[21741];
assign MEM[39165] = MEM[21738] + MEM[21858];
assign MEM[39166] = MEM[21739] + MEM[21860];
assign MEM[39167] = MEM[21740] + MEM[21827];
assign MEM[39168] = MEM[21744] + MEM[21760];
assign MEM[39169] = MEM[21748] + MEM[21826];
assign MEM[39170] = MEM[21749] + MEM[21772];
assign MEM[39171] = MEM[21750] + MEM[21754];
assign MEM[39172] = MEM[21752] + MEM[21809];
assign MEM[39173] = MEM[21753] + MEM[21848];
assign MEM[39174] = MEM[21761] + MEM[21822];
assign MEM[39175] = MEM[21767] + MEM[21965];
assign MEM[39176] = MEM[21769] + MEM[21840];
assign MEM[39177] = MEM[21770] + MEM[21872];
assign MEM[39178] = MEM[21771] + MEM[21885];
assign MEM[39179] = MEM[21773] + MEM[21791];
assign MEM[39180] = MEM[21776] + MEM[21878];
assign MEM[39181] = MEM[21777] + MEM[21959];
assign MEM[39182] = MEM[21780] + MEM[21805];
assign MEM[39183] = MEM[21781] + MEM[21788];
assign MEM[39184] = MEM[21782] + MEM[21818];
assign MEM[39185] = MEM[21783] + MEM[21784];
assign MEM[39186] = MEM[21785] + MEM[21847];
assign MEM[39187] = MEM[21792] + MEM[21819];
assign MEM[39188] = MEM[21793] + MEM[21951];
assign MEM[39189] = MEM[21796] + MEM[21890];
assign MEM[39190] = MEM[21797] + MEM[21868];
assign MEM[39191] = MEM[21799] + MEM[21821];
assign MEM[39192] = MEM[21800] + MEM[21887];
assign MEM[39193] = MEM[21804] + MEM[21940];
assign MEM[39194] = MEM[21808] + MEM[21880];
assign MEM[39195] = MEM[21810] + MEM[21813];
assign MEM[39196] = MEM[21811] + MEM[21839];
assign MEM[39197] = MEM[21814] + MEM[21870];
assign MEM[39198] = MEM[21815] + MEM[21888];
assign MEM[39199] = MEM[21816] + MEM[22014];
assign MEM[39200] = MEM[21820] + MEM[21942];
assign MEM[39201] = MEM[21823] + MEM[21824];
assign MEM[39202] = MEM[21828] + MEM[21863];
assign MEM[39203] = MEM[21830] + MEM[22083];
assign MEM[39204] = MEM[21831] + MEM[22039];
assign MEM[39205] = MEM[21833] + MEM[21844];
assign MEM[39206] = MEM[21834] + MEM[22011];
assign MEM[39207] = MEM[21835] + MEM[21964];
assign MEM[39208] = MEM[21837] + MEM[21842];
assign MEM[39209] = MEM[21838] + MEM[21849];
assign MEM[39210] = MEM[21843] + MEM[21919];
assign MEM[39211] = MEM[21845] + MEM[21853];
assign MEM[39212] = MEM[21850] + MEM[21911];
assign MEM[39213] = MEM[21851] + MEM[21873];
assign MEM[39214] = MEM[21852] + MEM[21896];
assign MEM[39215] = MEM[21855] + MEM[21864];
assign MEM[39216] = MEM[21857] + MEM[21897];
assign MEM[39217] = MEM[21859] + MEM[21917];
assign MEM[39218] = MEM[21861] + MEM[21949];
assign MEM[39219] = MEM[21865] + MEM[21907];
assign MEM[39220] = MEM[21866] + MEM[22002];
assign MEM[39221] = MEM[21869] + MEM[21877];
assign MEM[39222] = MEM[21874] + MEM[21876];
assign MEM[39223] = MEM[21879] + MEM[21928];
assign MEM[39224] = MEM[21881] + MEM[21915];
assign MEM[39225] = MEM[21882] + MEM[22133];
assign MEM[39226] = MEM[21883] + MEM[21983];
assign MEM[39227] = MEM[21884] + MEM[21946];
assign MEM[39228] = MEM[21889] + MEM[21929];
assign MEM[39229] = MEM[21892] + MEM[21993];
assign MEM[39230] = MEM[21893] + MEM[21923];
assign MEM[39231] = MEM[21898] + MEM[22068];
assign MEM[39232] = MEM[21899] + MEM[21930];
assign MEM[39233] = MEM[21900] + MEM[22120];
assign MEM[39234] = MEM[21901] + MEM[21913];
assign MEM[39235] = MEM[21902] + MEM[21921];
assign MEM[39236] = MEM[21903] + MEM[21996];
assign MEM[39237] = MEM[21904] + MEM[21922];
assign MEM[39238] = MEM[21905] + MEM[21987];
assign MEM[39239] = MEM[21908] + MEM[21938];
assign MEM[39240] = MEM[21912] + MEM[22147];
assign MEM[39241] = MEM[21914] + MEM[21945];
assign MEM[39242] = MEM[21916] + MEM[21994];
assign MEM[39243] = MEM[21918] + MEM[21947];
assign MEM[39244] = MEM[21931] + MEM[21981];
assign MEM[39245] = MEM[21932] + MEM[21933];
assign MEM[39246] = MEM[21935] + MEM[21976];
assign MEM[39247] = MEM[21936] + MEM[22079];
assign MEM[39248] = MEM[21937] + MEM[21967];
assign MEM[39249] = MEM[21941] + MEM[22104];
assign MEM[39250] = MEM[21943] + MEM[21974];
assign MEM[39251] = MEM[21944] + MEM[21995];
assign MEM[39252] = MEM[21948] + MEM[22096];
assign MEM[39253] = MEM[21950] + MEM[21952];
assign MEM[39254] = MEM[21953] + MEM[22163];
assign MEM[39255] = MEM[21954] + MEM[21960];
assign MEM[39256] = MEM[21956] + MEM[22127];
assign MEM[39257] = MEM[21957] + MEM[21997];
assign MEM[39258] = MEM[21961] + MEM[22153];
assign MEM[39259] = MEM[21962] + MEM[21966];
assign MEM[39260] = MEM[21963] + MEM[22122];
assign MEM[39261] = MEM[21968] + MEM[21990];
assign MEM[39262] = MEM[21969] + MEM[22020];
assign MEM[39263] = MEM[21972] + MEM[21986];
assign MEM[39264] = MEM[21973] + MEM[22042];
assign MEM[39265] = MEM[21975] + MEM[22038];
assign MEM[39266] = MEM[21978] + MEM[22026];
assign MEM[39267] = MEM[21979] + MEM[22030];
assign MEM[39268] = MEM[21982] + MEM[22072];
assign MEM[39269] = MEM[21984] + MEM[22094];
assign MEM[39270] = MEM[21985] + MEM[22007];
assign MEM[39271] = MEM[21988] + MEM[22031];
assign MEM[39272] = MEM[21991] + MEM[22025];
assign MEM[39273] = MEM[21992] + MEM[22069];
assign MEM[39274] = MEM[21998] + MEM[22177];
assign MEM[39275] = MEM[21999] + MEM[22006];
assign MEM[39276] = MEM[22001] + MEM[22024];
assign MEM[39277] = MEM[22004] + MEM[22089];
assign MEM[39278] = MEM[22005] + MEM[22047];
assign MEM[39279] = MEM[22009] + MEM[22126];
assign MEM[39280] = MEM[22010] + MEM[22049];
assign MEM[39281] = MEM[22015] + MEM[22167];
assign MEM[39282] = MEM[22017] + MEM[22086];
assign MEM[39283] = MEM[22018] + MEM[22073];
assign MEM[39284] = MEM[22021] + MEM[22027];
assign MEM[39285] = MEM[22022] + MEM[22046];
assign MEM[39286] = MEM[22028] + MEM[22164];
assign MEM[39287] = MEM[22029] + MEM[22211];
assign MEM[39288] = MEM[22035] + MEM[22065];
assign MEM[39289] = MEM[22036] + MEM[22100];
assign MEM[39290] = MEM[22037] + MEM[22074];
assign MEM[39291] = MEM[22040] + MEM[22245];
assign MEM[39292] = MEM[22041] + MEM[22045];
assign MEM[39293] = MEM[22043] + MEM[22063];
assign MEM[39294] = MEM[22044] + MEM[22259];
assign MEM[39295] = MEM[22048] + MEM[22098];
assign MEM[39296] = MEM[22050] + MEM[22108];
assign MEM[39297] = MEM[22051] + MEM[22053];
assign MEM[39298] = MEM[22052] + MEM[22067];
assign MEM[39299] = MEM[22054] + MEM[22066];
assign MEM[39300] = MEM[22055] + MEM[22208];
assign MEM[39301] = MEM[22056] + MEM[22091];
assign MEM[39302] = MEM[22057] + MEM[22080];
assign MEM[39303] = MEM[22058] + MEM[22156];
assign MEM[39304] = MEM[22059] + MEM[22200];
assign MEM[39305] = MEM[22060] + MEM[22076];
assign MEM[39306] = MEM[22061] + MEM[22070];
assign MEM[39307] = MEM[22062] + MEM[22093];
assign MEM[39308] = MEM[22064] + MEM[22132];
assign MEM[39309] = MEM[22071] + MEM[22099];
assign MEM[39310] = MEM[22075] + MEM[22124];
assign MEM[39311] = MEM[22077] + MEM[22158];
assign MEM[39312] = MEM[22078] + MEM[22095];
assign MEM[39313] = MEM[22081] + MEM[22140];
assign MEM[39314] = MEM[22082] + MEM[22090];
assign MEM[39315] = MEM[22085] + MEM[22185];
assign MEM[39316] = MEM[22087] + MEM[22188];
assign MEM[39317] = MEM[22088] + MEM[22135];
assign MEM[39318] = MEM[22092] + MEM[22106];
assign MEM[39319] = MEM[22101] + MEM[22168];
assign MEM[39320] = MEM[22102] + MEM[22103];
assign MEM[39321] = MEM[22105] + MEM[22116];
assign MEM[39322] = MEM[22107] + MEM[22174];
assign MEM[39323] = MEM[22109] + MEM[22121];
assign MEM[39324] = MEM[22111] + MEM[22178];
assign MEM[39325] = MEM[22113] + MEM[22350];
assign MEM[39326] = MEM[22114] + MEM[22128];
assign MEM[39327] = MEM[22115] + MEM[22269];
assign MEM[39328] = MEM[22117] + MEM[22180];
assign MEM[39329] = MEM[22123] + MEM[22215];
assign MEM[39330] = MEM[22125] + MEM[22220];
assign MEM[39331] = MEM[22129] + MEM[22318];
assign MEM[39332] = MEM[22130] + MEM[22161];
assign MEM[39333] = MEM[22134] + MEM[22197];
assign MEM[39334] = MEM[22136] + MEM[22298];
assign MEM[39335] = MEM[22137] + MEM[22169];
assign MEM[39336] = MEM[22138] + MEM[22279];
assign MEM[39337] = MEM[22139] + MEM[22421];
assign MEM[39338] = MEM[22141] + MEM[22152];
assign MEM[39339] = MEM[22143] + MEM[22165];
assign MEM[39340] = MEM[22144] + MEM[22186];
assign MEM[39341] = MEM[22145] + MEM[22160];
assign MEM[39342] = MEM[22146] + MEM[22236];
assign MEM[39343] = MEM[22151] + MEM[22294];
assign MEM[39344] = MEM[22154] + MEM[22182];
assign MEM[39345] = MEM[22155] + MEM[22157];
assign MEM[39346] = MEM[22159] + MEM[22192];
assign MEM[39347] = MEM[22162] + MEM[22171];
assign MEM[39348] = MEM[22166] + MEM[22527];
assign MEM[39349] = MEM[22172] + MEM[22173];
assign MEM[39350] = MEM[22175] + MEM[22207];
assign MEM[39351] = MEM[22176] + MEM[22312];
assign MEM[39352] = MEM[22179] + MEM[22189];
assign MEM[39353] = MEM[22183] + MEM[22205];
assign MEM[39354] = MEM[22187] + MEM[22191];
assign MEM[39355] = MEM[22190] + MEM[22272];
assign MEM[39356] = MEM[22193] + MEM[22339];
assign MEM[39357] = MEM[22194] + MEM[22590];
assign MEM[39358] = MEM[22195] + MEM[22297];
assign MEM[39359] = MEM[22198] + MEM[22253];
assign MEM[39360] = MEM[22201] + MEM[22270];
assign MEM[39361] = MEM[22202] + MEM[22217];
assign MEM[39362] = MEM[22204] + MEM[22233];
assign MEM[39363] = MEM[22206] + MEM[22387];
assign MEM[39364] = MEM[22209] + MEM[22314];
assign MEM[39365] = MEM[22210] + MEM[22221];
assign MEM[39366] = MEM[22212] + MEM[22290];
assign MEM[39367] = MEM[22213] + MEM[22321];
assign MEM[39368] = MEM[22214] + MEM[22437];
assign MEM[39369] = MEM[22216] + MEM[22306];
assign MEM[39370] = MEM[22218] + MEM[22302];
assign MEM[39371] = MEM[22219] + MEM[22246];
assign MEM[39372] = MEM[22222] + MEM[22251];
assign MEM[39373] = MEM[22223] + MEM[22232];
assign MEM[39374] = MEM[22224] + MEM[22230];
assign MEM[39375] = MEM[22225] + MEM[22228];
assign MEM[39376] = MEM[22226] + MEM[22234];
assign MEM[39377] = MEM[22235] + MEM[22408];
assign MEM[39378] = MEM[22237] + MEM[22274];
assign MEM[39379] = MEM[22239] + MEM[22330];
assign MEM[39380] = MEM[22240] + MEM[22263];
assign MEM[39381] = MEM[22241] + MEM[22289];
assign MEM[39382] = MEM[22242] + MEM[22252];
assign MEM[39383] = MEM[22243] + MEM[22311];
assign MEM[39384] = MEM[22244] + MEM[22355];
assign MEM[39385] = MEM[22247] + MEM[22400];
assign MEM[39386] = MEM[22248] + MEM[22329];
assign MEM[39387] = MEM[22249] + MEM[22284];
assign MEM[39388] = MEM[22250] + MEM[22280];
assign MEM[39389] = MEM[22254] + MEM[22261];
assign MEM[39390] = MEM[22255] + MEM[22303];
assign MEM[39391] = MEM[22256] + MEM[22304];
assign MEM[39392] = MEM[22257] + MEM[22319];
assign MEM[39393] = MEM[22260] + MEM[22388];
assign MEM[39394] = MEM[22262] + MEM[22323];
assign MEM[39395] = MEM[22265] + MEM[22370];
assign MEM[39396] = MEM[22266] + MEM[22273];
assign MEM[39397] = MEM[22267] + MEM[22320];
assign MEM[39398] = MEM[22271] + MEM[22299];
assign MEM[39399] = MEM[22275] + MEM[22336];
assign MEM[39400] = MEM[22276] + MEM[22296];
assign MEM[39401] = MEM[22277] + MEM[22352];
assign MEM[39402] = MEM[22278] + MEM[22386];
assign MEM[39403] = MEM[22281] + MEM[22353];
assign MEM[39404] = MEM[22282] + MEM[22479];
assign MEM[39405] = MEM[22285] + MEM[22529];
assign MEM[39406] = MEM[22286] + MEM[22337];
assign MEM[39407] = MEM[22287] + MEM[22331];
assign MEM[39408] = MEM[22291] + MEM[22308];
assign MEM[39409] = MEM[22292] + MEM[22430];
assign MEM[39410] = MEM[22301] + MEM[22508];
assign MEM[39411] = MEM[22305] + MEM[22409];
assign MEM[39412] = MEM[22307] + MEM[22325];
assign MEM[39413] = MEM[22309] + MEM[22579];
assign MEM[39414] = MEM[22310] + MEM[22363];
assign MEM[39415] = MEM[22315] + MEM[22346];
assign MEM[39416] = MEM[22316] + MEM[22436];
assign MEM[39417] = MEM[22322] + MEM[22389];
assign MEM[39418] = MEM[22324] + MEM[22359];
assign MEM[39419] = MEM[22326] + MEM[22342];
assign MEM[39420] = MEM[22328] + MEM[22361];
assign MEM[39421] = MEM[22332] + MEM[22469];
assign MEM[39422] = MEM[22333] + MEM[22356];
assign MEM[39423] = MEM[22334] + MEM[22432];
assign MEM[39424] = MEM[22335] + MEM[22535];
assign MEM[39425] = MEM[22338] + MEM[22383];
assign MEM[39426] = MEM[22340] + MEM[22402];
assign MEM[39427] = MEM[22343] + MEM[22396];
assign MEM[39428] = MEM[22344] + MEM[22395];
assign MEM[39429] = MEM[22347] + MEM[22593];
assign MEM[39430] = MEM[22348] + MEM[22375];
assign MEM[39431] = MEM[22351] + MEM[22450];
assign MEM[39432] = MEM[22354] + MEM[22413];
assign MEM[39433] = MEM[22358] + MEM[22362];
assign MEM[39434] = MEM[22360] + MEM[22443];
assign MEM[39435] = MEM[22364] + MEM[22371];
assign MEM[39436] = MEM[22365] + MEM[22403];
assign MEM[39437] = MEM[22366] + MEM[22381];
assign MEM[39438] = MEM[22367] + MEM[22412];
assign MEM[39439] = MEM[22372] + MEM[22785];
assign MEM[39440] = MEM[22373] + MEM[22380];
assign MEM[39441] = MEM[22376] + MEM[22415];
assign MEM[39442] = MEM[22377] + MEM[22391];
assign MEM[39443] = MEM[22378] + MEM[22379];
assign MEM[39444] = MEM[22382] + MEM[22406];
assign MEM[39445] = MEM[22384] + MEM[22424];
assign MEM[39446] = MEM[22385] + MEM[22422];
assign MEM[39447] = MEM[22390] + MEM[22478];
assign MEM[39448] = MEM[22392] + MEM[22411];
assign MEM[39449] = MEM[22393] + MEM[22545];
assign MEM[39450] = MEM[22394] + MEM[22465];
assign MEM[39451] = MEM[22397] + MEM[22484];
assign MEM[39452] = MEM[22399] + MEM[22481];
assign MEM[39453] = MEM[22401] + MEM[22435];
assign MEM[39454] = MEM[22404] + MEM[22520];
assign MEM[39455] = MEM[22405] + MEM[22444];
assign MEM[39456] = MEM[22410] + MEM[22648];
assign MEM[39457] = MEM[22414] + MEM[22566];
assign MEM[39458] = MEM[22416] + MEM[22472];
assign MEM[39459] = MEM[22418] + MEM[22451];
assign MEM[39460] = MEM[22423] + MEM[22502];
assign MEM[39461] = MEM[22426] + MEM[22433];
assign MEM[39462] = MEM[22427] + MEM[22457];
assign MEM[39463] = MEM[22428] + MEM[22445];
assign MEM[39464] = MEM[22429] + MEM[22487];
assign MEM[39465] = MEM[22431] + MEM[22441];
assign MEM[39466] = MEM[22434] + MEM[22496];
assign MEM[39467] = MEM[22439] + MEM[22495];
assign MEM[39468] = MEM[22440] + MEM[22622];
assign MEM[39469] = MEM[22447] + MEM[22456];
assign MEM[39470] = MEM[22448] + MEM[22555];
assign MEM[39471] = MEM[22452] + MEM[22490];
assign MEM[39472] = MEM[22453] + MEM[22526];
assign MEM[39473] = MEM[22454] + MEM[22462];
assign MEM[39474] = MEM[22455] + MEM[22461];
assign MEM[39475] = MEM[22458] + MEM[22500];
assign MEM[39476] = MEM[22459] + MEM[22596];
assign MEM[39477] = MEM[22460] + MEM[22549];
assign MEM[39478] = MEM[22463] + MEM[22476];
assign MEM[39479] = MEM[22464] + MEM[22608];
assign MEM[39480] = MEM[22466] + MEM[22467];
assign MEM[39481] = MEM[22470] + MEM[22857];
assign MEM[39482] = MEM[22471] + MEM[22503];
assign MEM[39483] = MEM[22473] + MEM[22513];
assign MEM[39484] = MEM[22474] + MEM[22530];
assign MEM[39485] = MEM[22477] + MEM[22603];
assign MEM[39486] = MEM[22480] + MEM[22587];
assign MEM[39487] = MEM[22482] + MEM[22489];
assign MEM[39488] = MEM[22483] + MEM[22634];
assign MEM[39489] = MEM[22485] + MEM[22524];
assign MEM[39490] = MEM[22486] + MEM[22516];
assign MEM[39491] = MEM[22488] + MEM[22492];
assign MEM[39492] = MEM[22491] + MEM[22504];
assign MEM[39493] = MEM[22493] + MEM[22533];
assign MEM[39494] = MEM[22494] + MEM[22505];
assign MEM[39495] = MEM[22497] + MEM[22729];
assign MEM[39496] = MEM[22498] + MEM[22567];
assign MEM[39497] = MEM[22499] + MEM[22506];
assign MEM[39498] = MEM[22501] + MEM[22554];
assign MEM[39499] = MEM[22507] + MEM[22673];
assign MEM[39500] = MEM[22512] + MEM[22572];
assign MEM[39501] = MEM[22517] + MEM[22694];
assign MEM[39502] = MEM[22518] + MEM[22638];
assign MEM[39503] = MEM[22519] + MEM[22557];
assign MEM[39504] = MEM[22521] + MEM[22645];
assign MEM[39505] = MEM[22522] + MEM[22525];
assign MEM[39506] = MEM[22523] + MEM[22556];
assign MEM[39507] = MEM[22528] + MEM[22541];
assign MEM[39508] = MEM[22531] + MEM[22551];
assign MEM[39509] = MEM[22532] + MEM[22646];
assign MEM[39510] = MEM[22534] + MEM[22546];
assign MEM[39511] = MEM[22536] + MEM[22605];
assign MEM[39512] = MEM[22537] + MEM[22606];
assign MEM[39513] = MEM[22538] + MEM[22571];
assign MEM[39514] = MEM[22539] + MEM[22620];
assign MEM[39515] = MEM[22540] + MEM[22624];
assign MEM[39516] = MEM[22542] + MEM[22650];
assign MEM[39517] = MEM[22543] + MEM[22568];
assign MEM[39518] = MEM[22544] + MEM[22599];
assign MEM[39519] = MEM[22547] + MEM[22621];
assign MEM[39520] = MEM[22548] + MEM[22756];
assign MEM[39521] = MEM[22550] + MEM[22662];
assign MEM[39522] = MEM[22558] + MEM[22601];
assign MEM[39523] = MEM[22559] + MEM[22615];
assign MEM[39524] = MEM[22560] + MEM[22693];
assign MEM[39525] = MEM[22561] + MEM[22618];
assign MEM[39526] = MEM[22563] + MEM[22602];
assign MEM[39527] = MEM[22565] + MEM[22631];
assign MEM[39528] = MEM[22570] + MEM[22688];
assign MEM[39529] = MEM[22573] + MEM[22611];
assign MEM[39530] = MEM[22574] + MEM[22765];
assign MEM[39531] = MEM[22577] + MEM[22644];
assign MEM[39532] = MEM[22578] + MEM[22589];
assign MEM[39533] = MEM[22581] + MEM[22755];
assign MEM[39534] = MEM[22582] + MEM[22751];
assign MEM[39535] = MEM[22583] + MEM[22668];
assign MEM[39536] = MEM[22584] + MEM[22667];
assign MEM[39537] = MEM[22585] + MEM[22659];
assign MEM[39538] = MEM[22588] + MEM[22690];
assign MEM[39539] = MEM[22591] + MEM[22640];
assign MEM[39540] = MEM[22592] + MEM[22808];
assign MEM[39541] = MEM[22594] + MEM[22666];
assign MEM[39542] = MEM[22595] + MEM[22636];
assign MEM[39543] = MEM[22597] + MEM[22691];
assign MEM[39544] = MEM[22598] + MEM[22701];
assign MEM[39545] = MEM[22604] + MEM[22671];
assign MEM[39546] = MEM[22607] + MEM[22616];
assign MEM[39547] = MEM[22609] + MEM[22763];
assign MEM[39548] = MEM[22610] + MEM[22613];
assign MEM[39549] = MEM[22612] + MEM[22750];
assign MEM[39550] = MEM[22614] + MEM[22875];
assign MEM[39551] = MEM[22619] + MEM[22989];
assign MEM[39552] = MEM[22626] + MEM[22647];
assign MEM[39553] = MEM[22628] + MEM[22700];
assign MEM[39554] = MEM[22629] + MEM[22637];
assign MEM[39555] = MEM[22630] + MEM[22641];
assign MEM[39556] = MEM[22632] + MEM[22856];
assign MEM[39557] = MEM[22635] + MEM[22780];
assign MEM[39558] = MEM[22639] + MEM[22669];
assign MEM[39559] = MEM[22643] + MEM[22884];
assign MEM[39560] = MEM[22649] + MEM[22682];
assign MEM[39561] = MEM[22653] + MEM[22657];
assign MEM[39562] = MEM[22654] + MEM[22722];
assign MEM[39563] = MEM[22656] + MEM[22664];
assign MEM[39564] = MEM[22658] + MEM[22786];
assign MEM[39565] = MEM[22660] + MEM[22723];
assign MEM[39566] = MEM[22663] + MEM[22705];
assign MEM[39567] = MEM[22672] + MEM[22708];
assign MEM[39568] = MEM[22674] + MEM[22846];
assign MEM[39569] = MEM[22675] + MEM[22861];
assign MEM[39570] = MEM[22676] + MEM[22807];
assign MEM[39571] = MEM[22677] + MEM[22895];
assign MEM[39572] = MEM[22678] + MEM[22679];
assign MEM[39573] = MEM[22681] + MEM[22799];
assign MEM[39574] = MEM[22683] + MEM[22684];
assign MEM[39575] = MEM[22685] + MEM[23005];
assign MEM[39576] = MEM[22686] + MEM[22689];
assign MEM[39577] = MEM[22687] + MEM[22706];
assign MEM[39578] = MEM[22695] + MEM[22744];
assign MEM[39579] = MEM[22696] + MEM[22871];
assign MEM[39580] = MEM[22697] + MEM[22698];
assign MEM[39581] = MEM[22699] + MEM[22711];
assign MEM[39582] = MEM[22704] + MEM[22716];
assign MEM[39583] = MEM[22707] + MEM[22880];
assign MEM[39584] = MEM[22712] + MEM[22735];
assign MEM[39585] = MEM[22714] + MEM[22896];
assign MEM[39586] = MEM[22715] + MEM[22802];
assign MEM[39587] = MEM[22717] + MEM[22939];
assign MEM[39588] = MEM[22718] + MEM[22732];
assign MEM[39589] = MEM[22719] + MEM[22782];
assign MEM[39590] = MEM[22720] + MEM[22770];
assign MEM[39591] = MEM[22724] + MEM[22795];
assign MEM[39592] = MEM[22726] + MEM[22862];
assign MEM[39593] = MEM[22727] + MEM[22743];
assign MEM[39594] = MEM[22728] + MEM[22813];
assign MEM[39595] = MEM[22731] + MEM[22737];
assign MEM[39596] = MEM[22733] + MEM[22734];
assign MEM[39597] = MEM[22738] + MEM[22742];
assign MEM[39598] = MEM[22739] + MEM[22815];
assign MEM[39599] = MEM[22740] + MEM[22800];
assign MEM[39600] = MEM[22745] + MEM[22776];
assign MEM[39601] = MEM[22747] + MEM[22778];
assign MEM[39602] = MEM[22748] + MEM[22760];
assign MEM[39603] = MEM[22749] + MEM[22752];
assign MEM[39604] = MEM[22753] + MEM[22775];
assign MEM[39605] = MEM[22754] + MEM[22814];
assign MEM[39606] = MEM[22757] + MEM[22843];
assign MEM[39607] = MEM[22758] + MEM[22830];
assign MEM[39608] = MEM[22759] + MEM[22764];
assign MEM[39609] = MEM[22767] + MEM[22818];
assign MEM[39610] = MEM[22768] + MEM[22824];
assign MEM[39611] = MEM[22769] + MEM[22771];
assign MEM[39612] = MEM[22773] + MEM[22899];
assign MEM[39613] = MEM[22774] + MEM[22866];
assign MEM[39614] = MEM[22777] + MEM[22801];
assign MEM[39615] = MEM[22779] + MEM[22832];
assign MEM[39616] = MEM[22781] + MEM[22834];
assign MEM[39617] = MEM[22783] + MEM[22852];
assign MEM[39618] = MEM[22787] + MEM[22793];
assign MEM[39619] = MEM[22788] + MEM[22845];
assign MEM[39620] = MEM[22789] + MEM[22819];
assign MEM[39621] = MEM[22790] + MEM[22831];
assign MEM[39622] = MEM[22791] + MEM[22933];
assign MEM[39623] = MEM[22792] + MEM[22833];
assign MEM[39624] = MEM[22794] + MEM[22806];
assign MEM[39625] = MEM[22796] + MEM[22964];
assign MEM[39626] = MEM[22797] + MEM[22878];
assign MEM[39627] = MEM[22798] + MEM[22817];
assign MEM[39628] = MEM[22803] + MEM[22859];
assign MEM[39629] = MEM[22804] + MEM[22838];
assign MEM[39630] = MEM[22805] + MEM[22836];
assign MEM[39631] = MEM[22809] + MEM[22898];
assign MEM[39632] = MEM[22810] + MEM[22886];
assign MEM[39633] = MEM[22811] + MEM[22863];
assign MEM[39634] = MEM[22812] + MEM[22820];
assign MEM[39635] = MEM[22816] + MEM[23147];
assign MEM[39636] = MEM[22821] + MEM[23086];
assign MEM[39637] = MEM[22822] + MEM[22868];
assign MEM[39638] = MEM[22823] + MEM[22867];
assign MEM[39639] = MEM[22825] + MEM[22931];
assign MEM[39640] = MEM[22826] + MEM[22855];
assign MEM[39641] = MEM[22827] + MEM[22842];
assign MEM[39642] = MEM[22828] + MEM[22925];
assign MEM[39643] = MEM[22829] + MEM[22839];
assign MEM[39644] = MEM[22837] + MEM[22887];
assign MEM[39645] = MEM[22840] + MEM[22848];
assign MEM[39646] = MEM[22841] + MEM[22954];
assign MEM[39647] = MEM[22844] + MEM[23003];
assign MEM[39648] = MEM[22847] + MEM[22949];
assign MEM[39649] = MEM[22850] + MEM[23130];
assign MEM[39650] = MEM[22851] + MEM[22998];
assign MEM[39651] = MEM[22853] + MEM[22858];
assign MEM[39652] = MEM[22854] + MEM[22870];
assign MEM[39653] = MEM[22860] + MEM[22986];
assign MEM[39654] = MEM[22864] + MEM[23057];
assign MEM[39655] = MEM[22865] + MEM[22872];
assign MEM[39656] = MEM[22873] + MEM[22915];
assign MEM[39657] = MEM[22874] + MEM[22904];
assign MEM[39658] = MEM[22876] + MEM[22914];
assign MEM[39659] = MEM[22877] + MEM[22885];
assign MEM[39660] = MEM[22879] + MEM[22909];
assign MEM[39661] = MEM[22881] + MEM[22968];
assign MEM[39662] = MEM[22882] + MEM[22918];
assign MEM[39663] = MEM[22888] + MEM[22936];
assign MEM[39664] = MEM[22889] + MEM[22922];
assign MEM[39665] = MEM[22890] + MEM[22908];
assign MEM[39666] = MEM[22891] + MEM[22913];
assign MEM[39667] = MEM[22892] + MEM[23075];
assign MEM[39668] = MEM[22893] + MEM[22953];
assign MEM[39669] = MEM[22894] + MEM[22919];
assign MEM[39670] = MEM[22897] + MEM[22970];
assign MEM[39671] = MEM[22900] + MEM[23009];
assign MEM[39672] = MEM[22901] + MEM[22912];
assign MEM[39673] = MEM[22902] + MEM[22928];
assign MEM[39674] = MEM[22903] + MEM[22958];
assign MEM[39675] = MEM[22905] + MEM[23013];
assign MEM[39676] = MEM[22906] + MEM[22910];
assign MEM[39677] = MEM[22907] + MEM[22940];
assign MEM[39678] = MEM[22911] + MEM[22963];
assign MEM[39679] = MEM[22916] + MEM[22947];
assign MEM[39680] = MEM[22917] + MEM[22965];
assign MEM[39681] = MEM[22920] + MEM[22935];
assign MEM[39682] = MEM[22921] + MEM[23105];
assign MEM[39683] = MEM[22923] + MEM[22966];
assign MEM[39684] = MEM[22924] + MEM[22962];
assign MEM[39685] = MEM[22926] + MEM[22990];
assign MEM[39686] = MEM[22927] + MEM[22948];
assign MEM[39687] = MEM[22929] + MEM[23015];
assign MEM[39688] = MEM[22930] + MEM[22952];
assign MEM[39689] = MEM[22932] + MEM[22994];
assign MEM[39690] = MEM[22934] + MEM[23016];
assign MEM[39691] = MEM[22937] + MEM[23029];
assign MEM[39692] = MEM[22938] + MEM[22979];
assign MEM[39693] = MEM[22941] + MEM[23074];
assign MEM[39694] = MEM[22942] + MEM[22960];
assign MEM[39695] = MEM[22943] + MEM[23050];
assign MEM[39696] = MEM[22944] + MEM[22951];
assign MEM[39697] = MEM[22945] + MEM[23096];
assign MEM[39698] = MEM[22946] + MEM[22974];
assign MEM[39699] = MEM[22950] + MEM[22997];
assign MEM[39700] = MEM[22955] + MEM[22959];
assign MEM[39701] = MEM[22956] + MEM[22972];
assign MEM[39702] = MEM[22957] + MEM[22984];
assign MEM[39703] = MEM[22961] + MEM[23165];
assign MEM[39704] = MEM[22967] + MEM[22971];
assign MEM[39705] = MEM[22969] + MEM[23066];
assign MEM[39706] = MEM[22973] + MEM[23174];
assign MEM[39707] = MEM[22975] + MEM[23253];
assign MEM[39708] = MEM[22976] + MEM[22985];
assign MEM[39709] = MEM[22977] + MEM[22992];
assign MEM[39710] = MEM[22978] + MEM[23000];
assign MEM[39711] = MEM[22980] + MEM[22982];
assign MEM[39712] = MEM[22981] + MEM[23036];
assign MEM[39713] = MEM[22983] + MEM[23014];
assign MEM[39714] = MEM[22987] + MEM[23087];
assign MEM[39715] = MEM[22988] + MEM[23001];
assign MEM[39716] = MEM[22991] + MEM[23031];
assign MEM[39717] = MEM[22993] + MEM[23025];
assign MEM[39718] = MEM[22995] + MEM[23004];
assign MEM[39719] = MEM[22996] + MEM[23020];
assign MEM[39720] = MEM[22999] + MEM[23019];
assign MEM[39721] = MEM[23002] + MEM[23044];
assign MEM[39722] = MEM[23006] + MEM[23187];
assign MEM[39723] = MEM[23007] + MEM[23038];
assign MEM[39724] = MEM[23008] + MEM[23052];
assign MEM[39725] = MEM[23010] + MEM[23135];
assign MEM[39726] = MEM[23011] + MEM[23055];
assign MEM[39727] = MEM[23012] + MEM[23073];
assign MEM[39728] = MEM[23017] + MEM[23030];
assign MEM[39729] = MEM[23018] + MEM[23202];
assign MEM[39730] = MEM[23021] + MEM[23035];
assign MEM[39731] = MEM[23022] + MEM[23079];
assign MEM[39732] = MEM[23023] + MEM[23034];
assign MEM[39733] = MEM[23024] + MEM[23027];
assign MEM[39734] = MEM[23026] + MEM[23058];
assign MEM[39735] = MEM[23028] + MEM[23041];
assign MEM[39736] = MEM[23032] + MEM[23113];
assign MEM[39737] = MEM[23033] + MEM[23039];
assign MEM[39738] = MEM[23037] + MEM[23069];
assign MEM[39739] = MEM[23040] + MEM[23047];
assign MEM[39740] = MEM[23042] + MEM[23319];
assign MEM[39741] = MEM[23043] + MEM[23053];
assign MEM[39742] = MEM[23045] + MEM[23062];
assign MEM[39743] = MEM[23046] + MEM[23241];
assign MEM[39744] = MEM[23048] + MEM[23095];
assign MEM[39745] = MEM[23049] + MEM[23094];
assign MEM[39746] = MEM[23051] + MEM[23091];
assign MEM[39747] = MEM[23054] + MEM[23078];
assign MEM[39748] = MEM[23056] + MEM[23080];
assign MEM[39749] = MEM[23059] + MEM[23123];
assign MEM[39750] = MEM[23060] + MEM[23136];
assign MEM[39751] = MEM[23061] + MEM[23077];
assign MEM[39752] = MEM[23063] + MEM[23100];
assign MEM[39753] = MEM[23064] + MEM[23082];
assign MEM[39754] = MEM[23065] + MEM[23104];
assign MEM[39755] = MEM[23067] + MEM[23286];
assign MEM[39756] = MEM[23068] + MEM[23220];
assign MEM[39757] = MEM[23070] + MEM[23155];
assign MEM[39758] = MEM[23071] + MEM[23122];
assign MEM[39759] = MEM[23072] + MEM[23081];
assign MEM[39760] = MEM[23076] + MEM[23180];
assign MEM[39761] = MEM[23083] + MEM[23084];
assign MEM[39762] = MEM[23085] + MEM[23153];
assign MEM[39763] = MEM[23088] + MEM[23146];
assign MEM[39764] = MEM[23089] + MEM[23128];
assign MEM[39765] = MEM[23090] + MEM[23168];
assign MEM[39766] = MEM[23092] + MEM[23199];
assign MEM[39767] = MEM[23093] + MEM[23342];
assign MEM[39768] = MEM[23097] + MEM[23161];
assign MEM[39769] = MEM[23098] + MEM[23109];
assign MEM[39770] = MEM[23099] + MEM[23246];
assign MEM[39771] = MEM[23101] + MEM[23178];
assign MEM[39772] = MEM[23102] + MEM[23203];
assign MEM[39773] = MEM[23103] + MEM[23185];
assign MEM[39774] = MEM[23106] + MEM[23114];
assign MEM[39775] = MEM[23107] + MEM[23196];
assign MEM[39776] = MEM[23108] + MEM[23317];
assign MEM[39777] = MEM[23110] + MEM[23217];
assign MEM[39778] = MEM[23111] + MEM[23173];
assign MEM[39779] = MEM[23112] + MEM[23195];
assign MEM[39780] = MEM[23115] + MEM[23133];
assign MEM[39781] = MEM[23116] + MEM[23142];
assign MEM[39782] = MEM[23117] + MEM[23149];
assign MEM[39783] = MEM[23118] + MEM[23137];
assign MEM[39784] = MEM[23119] + MEM[23172];
assign MEM[39785] = MEM[23120] + MEM[23129];
assign MEM[39786] = MEM[23121] + MEM[23131];
assign MEM[39787] = MEM[23124] + MEM[23132];
assign MEM[39788] = MEM[23125] + MEM[23154];
assign MEM[39789] = MEM[23126] + MEM[23248];
assign MEM[39790] = MEM[23127] + MEM[23143];
assign MEM[39791] = MEM[23134] + MEM[23157];
assign MEM[39792] = MEM[23138] + MEM[23156];
assign MEM[39793] = MEM[23139] + MEM[23158];
assign MEM[39794] = MEM[23140] + MEM[23236];
assign MEM[39795] = MEM[23141] + MEM[23183];
assign MEM[39796] = MEM[23144] + MEM[23225];
assign MEM[39797] = MEM[23145] + MEM[23151];
assign MEM[39798] = MEM[23148] + MEM[23177];
assign MEM[39799] = MEM[23150] + MEM[23167];
assign MEM[39800] = MEM[23152] + MEM[23182];
assign MEM[39801] = MEM[23159] + MEM[23192];
assign MEM[39802] = MEM[23160] + MEM[23219];
assign MEM[39803] = MEM[23162] + MEM[23169];
assign MEM[39804] = MEM[23163] + MEM[23218];
assign MEM[39805] = MEM[23164] + MEM[23237];
assign MEM[39806] = MEM[23166] + MEM[23232];
assign MEM[39807] = MEM[23170] + MEM[23228];
assign MEM[39808] = MEM[23171] + MEM[23181];
assign MEM[39809] = MEM[23175] + MEM[24336];
assign MEM[39810] = MEM[23176] + MEM[23207];
assign MEM[39811] = MEM[23179] + MEM[23189];
assign MEM[39812] = MEM[23184] + MEM[23194];
assign MEM[39813] = MEM[23186] + MEM[23211];
assign MEM[39814] = MEM[23188] + MEM[23201];
assign MEM[39815] = MEM[23190] + MEM[23366];
assign MEM[39816] = MEM[23191] + MEM[23298];
assign MEM[39817] = MEM[23193] + MEM[23255];
assign MEM[39818] = MEM[23197] + MEM[23335];
assign MEM[39819] = MEM[23198] + MEM[23280];
assign MEM[39820] = MEM[23200] + MEM[23233];
assign MEM[39821] = MEM[23204] + MEM[23278];
assign MEM[39822] = MEM[23205] + MEM[23222];
assign MEM[39823] = MEM[23206] + MEM[23333];
assign MEM[39824] = MEM[23208] + MEM[26491];
assign MEM[39825] = MEM[23209] + MEM[23829];
assign MEM[39826] = MEM[23210] + MEM[23284];
assign MEM[39827] = MEM[23212] + MEM[23239];
assign MEM[39828] = MEM[23213] + MEM[23265];
assign MEM[39829] = MEM[23214] + MEM[23215];
assign MEM[39830] = MEM[23216] + MEM[23289];
assign MEM[39831] = MEM[23221] + MEM[23997];
assign MEM[39832] = MEM[23223] + MEM[23964];
assign MEM[39833] = MEM[23224] + MEM[23273];
assign MEM[39834] = MEM[23226] + MEM[23279];
assign MEM[39835] = MEM[23227] + MEM[23251];
assign MEM[39836] = MEM[23229] + MEM[23293];
assign MEM[39837] = MEM[23230] + MEM[23272];
assign MEM[39838] = MEM[23231] + MEM[23297];
assign MEM[39839] = MEM[23234] + MEM[23247];
assign MEM[39840] = MEM[23235] + MEM[23244];
assign MEM[39841] = MEM[23238] + MEM[27562];
assign MEM[39842] = MEM[23240] + MEM[23274];
assign MEM[39843] = MEM[23242] + MEM[23259];
assign MEM[39844] = MEM[23245] + MEM[23287];
assign MEM[39845] = MEM[23249] + MEM[23558];
assign MEM[39846] = MEM[23250] + MEM[23305];
assign MEM[39847] = MEM[23252] + MEM[24910];
assign MEM[39848] = MEM[23254] + MEM[23268];
assign MEM[39849] = MEM[23256] + MEM[23269];
assign MEM[39850] = MEM[23257] + MEM[23314];
assign MEM[39851] = MEM[23258] + MEM[23260];
assign MEM[39852] = MEM[23261] + MEM[23343];
assign MEM[39853] = MEM[23262] + MEM[23267];
assign MEM[39854] = MEM[23263] + MEM[23266];
assign MEM[39855] = MEM[23264] + MEM[23307];
assign MEM[39856] = MEM[23270] + MEM[23347];
assign MEM[39857] = MEM[23271] + MEM[23316];
assign MEM[39858] = MEM[23275] + MEM[24114];
assign MEM[39859] = MEM[23276] + MEM[23285];
assign MEM[39860] = MEM[23277] + MEM[23900];
assign MEM[39861] = MEM[23281] + MEM[23889];
assign MEM[39862] = MEM[23282] + MEM[23315];
assign MEM[39863] = MEM[23283] + MEM[23364];
assign MEM[39864] = MEM[23288] + MEM[23300];
assign MEM[39865] = MEM[23290] + MEM[23338];
assign MEM[39866] = MEM[23291] + MEM[26572];
assign MEM[39867] = MEM[23292] + MEM[23294];
assign MEM[39868] = MEM[23295] + MEM[23685];
assign MEM[39869] = MEM[23296] + MEM[23336];
assign MEM[39870] = MEM[23299] + MEM[23805];
assign MEM[39871] = MEM[23301] + MEM[23304];
assign MEM[39872] = MEM[23302] + MEM[23329];
assign MEM[39873] = MEM[23303] + MEM[23659];
assign MEM[39874] = MEM[23306] + MEM[23310];
assign MEM[39875] = MEM[23308] + MEM[23359];
assign MEM[39876] = MEM[23309] + MEM[23325];
assign MEM[39877] = MEM[23311] + MEM[23340];
assign MEM[39878] = MEM[23312] + MEM[23351];
assign MEM[39879] = MEM[23313] + MEM[23902];
assign MEM[39880] = MEM[23318] + MEM[23940];
assign MEM[39881] = MEM[23320] + MEM[23355];
assign MEM[39882] = MEM[23321] + MEM[24921];
assign MEM[39883] = MEM[23322] + MEM[23354];
assign MEM[39884] = MEM[23323] + MEM[23353];
assign MEM[39885] = MEM[23324] + MEM[23332];
assign MEM[39886] = MEM[23326] + MEM[23339];
assign MEM[39887] = MEM[23327] + MEM[23360];
assign MEM[39888] = MEM[23328] + MEM[24892];
assign MEM[39889] = MEM[23330] + MEM[23334];
assign MEM[39890] = MEM[23331] + MEM[24001];
assign MEM[39891] = MEM[23337] + MEM[23805];
assign MEM[39892] = MEM[23341] + MEM[24180];
assign MEM[39893] = MEM[23344] + MEM[24146];
assign MEM[39894] = MEM[23345] + MEM[24120];
assign MEM[39895] = MEM[23346] + MEM[23684];
assign MEM[39896] = MEM[23348] + MEM[26239];
assign MEM[39897] = MEM[23349] + MEM[24001];
assign MEM[39898] = MEM[23350] + MEM[24280];
assign MEM[39899] = MEM[23352] + MEM[23358];
assign MEM[39900] = MEM[23356] + MEM[24146];
assign MEM[39901] = MEM[23357] + MEM[25578];
assign MEM[39902] = MEM[23361] + MEM[24700];
assign MEM[39903] = MEM[23362] + MEM[23888];
assign MEM[39904] = MEM[23363] + MEM[23829];
assign MEM[39905] = MEM[23366] + MEM[25398];
assign MEM[39906] = MEM[23391] + MEM[24082];
assign MEM[39907] = MEM[23391] + MEM[24328];
assign MEM[39908] = MEM[23430] + MEM[23964];
assign MEM[39909] = MEM[23430] + MEM[25318];
assign MEM[39910] = MEM[23487] + MEM[24485];
assign MEM[39911] = MEM[23487] + MEM[25849];
assign MEM[39912] = MEM[23558] + MEM[23889];
assign MEM[39913] = MEM[23659] + MEM[23759];
assign MEM[39914] = MEM[23684] + MEM[25854];
assign MEM[39915] = MEM[23685] + MEM[25178];
assign MEM[39916] = MEM[23759] + MEM[24120];
assign MEM[39917] = MEM[23888] + MEM[23891];
assign MEM[39918] = MEM[23891] + MEM[26176];
assign MEM[39919] = MEM[23900] + MEM[25178];
assign MEM[39920] = MEM[23902] + MEM[24180];
assign MEM[39921] = MEM[23940] + MEM[24160];
assign MEM[39922] = MEM[23997] + MEM[25398];
assign MEM[39923] = MEM[24082] + MEM[24211];
assign MEM[39924] = MEM[24085] + MEM[24356];
assign MEM[39925] = MEM[24085] + MEM[26722];
assign MEM[39926] = MEM[24095] + MEM[26015];
assign MEM[39927] = MEM[24095] + MEM[26677];
assign MEM[39928] = MEM[24114] + MEM[24830];
assign MEM[39929] = MEM[24160] + MEM[24643];
assign MEM[39930] = MEM[24167] + MEM[24204];
assign MEM[39931] = MEM[24167] + MEM[24780];
assign MEM[39932] = MEM[24179] + MEM[24189];
assign MEM[39933] = MEM[24179] + MEM[24212];
assign MEM[39934] = MEM[24189] + MEM[24700];
assign MEM[39935] = MEM[24204] + MEM[24981];
assign MEM[39936] = MEM[24211] + MEM[24605];
assign MEM[39937] = MEM[24212] + MEM[24280];
assign MEM[39938] = MEM[24297] + MEM[24849];
assign MEM[39939] = MEM[24297] + MEM[24981];
assign MEM[39940] = MEM[24328] + MEM[25909];
assign MEM[39941] = MEM[24336] + MEM[24815];
assign MEM[39942] = MEM[24356] + MEM[24747];
assign MEM[39943] = MEM[24394] + MEM[24449];
assign MEM[39944] = MEM[24394] + MEM[25476];
assign MEM[39945] = MEM[24449] + MEM[24540];
assign MEM[39946] = MEM[24485] + MEM[24747];
assign MEM[39947] = MEM[24540] + MEM[26171];
assign MEM[39948] = MEM[24600] + MEM[24756];
assign MEM[39949] = MEM[24600] + MEM[26587];
assign MEM[39950] = MEM[24605] + MEM[29829];
assign MEM[39951] = MEM[24643] + MEM[27055];
assign MEM[39952] = MEM[24718] + MEM[25285];
assign MEM[39953] = MEM[24718] + MEM[25635];
assign MEM[39954] = MEM[24756] + MEM[26801];
assign MEM[39955] = MEM[24780] + MEM[26407];
assign MEM[39956] = MEM[24815] + MEM[24830];
assign MEM[39957] = MEM[24849] + MEM[28683];
assign MEM[39958] = MEM[24851] + MEM[25635];
assign MEM[39959] = MEM[24851] + MEM[25723];
assign MEM[39960] = MEM[24892] + MEM[26157];
assign MEM[39961] = MEM[24910] + MEM[25581];
assign MEM[39962] = MEM[24921] + MEM[28191];
assign MEM[39963] = MEM[24964] + MEM[25230];
assign MEM[39964] = MEM[24964] + MEM[25285];
assign MEM[39965] = MEM[24997] + MEM[25523];
assign MEM[39966] = MEM[24997] + MEM[25855];
assign MEM[39967] = MEM[25230] + MEM[25909];
assign MEM[39968] = MEM[25263] + MEM[25709];
assign MEM[39969] = MEM[25263] + MEM[26077];
assign MEM[39970] = MEM[25266] + MEM[27087];
assign MEM[39971] = MEM[25266] + MEM[27452];
assign MEM[39972] = MEM[25318] + MEM[25628];
assign MEM[39973] = MEM[25327] + MEM[25581];
assign MEM[39974] = MEM[25327] + MEM[26328];
assign MEM[39975] = MEM[25367] + MEM[25855];
assign MEM[39976] = MEM[25367] + MEM[26156];
assign MEM[39977] = MEM[25444] + MEM[26048];
assign MEM[39978] = MEM[25444] + MEM[26382];
assign MEM[39979] = MEM[25476] + MEM[26271];
assign MEM[39980] = MEM[25481] + MEM[25863];
assign MEM[39981] = MEM[25481] + MEM[27007];
assign MEM[39982] = MEM[25523] + MEM[25578];
assign MEM[39983] = MEM[25628] + MEM[26293];
assign MEM[39984] = MEM[25709] + MEM[26015];
assign MEM[39985] = MEM[25723] + MEM[26897];
assign MEM[39986] = MEM[25849] + MEM[26798];
assign MEM[39987] = MEM[25854] + MEM[26417];
assign MEM[39988] = MEM[25863] + MEM[26391];
assign MEM[39989] = MEM[26020] + MEM[26157];
assign MEM[39990] = MEM[26020] + MEM[27310];
assign MEM[39991] = MEM[26040] + MEM[26310];
assign MEM[39992] = MEM[26040] + MEM[28344];
assign MEM[39993] = MEM[26048] + MEM[26901];
assign MEM[39994] = MEM[26077] + MEM[26312];
assign MEM[39995] = MEM[26156] + MEM[26246];
assign MEM[39996] = MEM[26171] + MEM[26677];
assign MEM[39997] = MEM[26176] + MEM[26716];
assign MEM[39998] = MEM[26192] + MEM[26239];
assign MEM[39999] = MEM[26192] + MEM[26410];
assign MEM[40000] = MEM[26194] + MEM[26328];
assign MEM[40001] = MEM[26194] + MEM[26789];
assign MEM[40002] = MEM[26205] + MEM[26587];
assign MEM[40003] = MEM[26205] + MEM[27110];
assign MEM[40004] = MEM[26207] + MEM[26259];
assign MEM[40005] = MEM[26207] + MEM[29793];
assign MEM[40006] = MEM[26246] + MEM[26483];
assign MEM[40007] = MEM[26259] + MEM[29841];
assign MEM[40008] = MEM[26271] + MEM[26644];
assign MEM[40009] = MEM[26293] + MEM[26547];
assign MEM[40010] = MEM[26310] + MEM[28555];
assign MEM[40011] = MEM[26312] + MEM[27310];
assign MEM[40012] = MEM[26335] + MEM[26461];
assign MEM[40013] = MEM[26335] + MEM[26491];
assign MEM[40014] = MEM[26382] + MEM[26798];
assign MEM[40015] = MEM[26391] + MEM[26740];
assign MEM[40016] = MEM[26407] + MEM[26897];
assign MEM[40017] = MEM[26410] + MEM[26461];
assign MEM[40018] = MEM[26417] + MEM[26686];
assign MEM[40019] = MEM[26483] + MEM[26788];
assign MEM[40020] = MEM[26547] + MEM[27022];
assign MEM[40021] = MEM[26572] + MEM[27024];
assign MEM[40022] = MEM[26611] + MEM[27265];
assign MEM[40023] = MEM[26611] + MEM[28466];
assign MEM[40024] = MEM[26644] + MEM[29748];
assign MEM[40025] = MEM[26650] + MEM[27022];
assign MEM[40026] = MEM[26650] + MEM[27303];
assign MEM[40027] = MEM[26686] + MEM[27173];
assign MEM[40028] = MEM[26716] + MEM[28524];
assign MEM[40029] = MEM[26722] + MEM[29175];
assign MEM[40030] = MEM[26740] + MEM[29639];
assign MEM[40031] = MEM[26788] + MEM[27240];
assign MEM[40032] = MEM[26789] + MEM[27335];
assign MEM[40033] = MEM[26801] + MEM[27125];
assign MEM[40034] = MEM[26901] + MEM[27110];
assign MEM[40035] = MEM[26903] + MEM[26934];
assign MEM[40036] = MEM[26903] + MEM[27329];
assign MEM[40037] = MEM[26934] + MEM[28360];
assign MEM[40038] = MEM[26964] + MEM[27007];
assign MEM[40039] = MEM[26964] + MEM[29784];
assign MEM[40040] = MEM[27024] + MEM[27249];
assign MEM[40041] = MEM[27055] + MEM[29531];
assign MEM[40042] = MEM[27083] + MEM[27303];
assign MEM[40043] = MEM[27083] + MEM[27452];
assign MEM[40044] = MEM[27087] + MEM[28021];
assign MEM[40045] = MEM[27118] + MEM[27154];
assign MEM[40046] = MEM[27118] + MEM[30019];
assign MEM[40047] = MEM[27125] + MEM[29553];
assign MEM[40048] = MEM[27152] + MEM[27173];
assign MEM[40049] = MEM[27152] + MEM[29312];
assign MEM[40050] = MEM[27154] + MEM[27669];
assign MEM[40051] = MEM[27240] + MEM[27588];
assign MEM[40052] = MEM[27249] + MEM[29368];
assign MEM[40053] = MEM[27265] + MEM[27559];
assign MEM[40054] = MEM[27329] + MEM[29801];
assign MEM[40055] = MEM[27335] + MEM[27447];
assign MEM[40056] = MEM[27447] + MEM[28933];
assign MEM[40057] = MEM[27559] + MEM[28979];
assign MEM[40058] = MEM[27562] + MEM[28344];
assign MEM[40059] = MEM[27588] + MEM[29086];
assign MEM[40060] = MEM[27650] + MEM[28499];
assign MEM[40061] = MEM[27650] + MEM[29312];
assign MEM[40062] = MEM[27669] + MEM[27826];
assign MEM[40063] = MEM[27826] + MEM[29773];
assign MEM[40064] = MEM[27949] + MEM[29134];
assign MEM[40065] = MEM[27949] + MEM[30093];
assign MEM[40066] = MEM[28021] + MEM[29086];
assign MEM[40067] = MEM[28191] + MEM[28466];
assign MEM[40068] = MEM[28230] + MEM[28555];
assign MEM[40069] = MEM[28230] + MEM[29885];
assign MEM[40070] = MEM[28293] + MEM[29347];
assign MEM[40071] = MEM[28293] + MEM[29788];
assign MEM[40072] = MEM[28360] + MEM[30061];
assign MEM[40073] = MEM[28499] + MEM[29750];
assign MEM[40074] = MEM[28504] + MEM[28803];
assign MEM[40075] = MEM[28504] + MEM[29480];
assign MEM[40076] = MEM[28524] + MEM[29811];
assign MEM[40077] = MEM[28683] + MEM[29271];
assign MEM[40078] = MEM[28738] + MEM[29368];
assign MEM[40079] = MEM[28738] + MEM[29722];
assign MEM[40080] = MEM[28803] + MEM[29745];
assign MEM[40081] = MEM[28910] + MEM[29713];
assign MEM[40082] = MEM[28910] + MEM[29982];
assign MEM[40083] = MEM[28933] + MEM[29763];
assign MEM[40084] = MEM[28979] + MEM[29244];
assign MEM[40085] = MEM[29121] + MEM[29271];
assign MEM[40086] = MEM[29121] + MEM[29708];
assign MEM[40087] = MEM[29134] + MEM[29780];
assign MEM[40088] = MEM[29175] + MEM[29932];
assign MEM[40089] = MEM[29241] + MEM[29347];
assign MEM[40090] = MEM[29241] + MEM[30065];
assign MEM[40091] = MEM[29244] + MEM[29435];
assign MEM[40092] = MEM[29325] + MEM[29694];
assign MEM[40093] = MEM[29325] + MEM[29748];
assign MEM[40094] = MEM[29410] + MEM[29733];
assign MEM[40095] = MEM[29410] + MEM[30093];
assign MEM[40096] = MEM[29435] + MEM[29847];
assign MEM[40097] = MEM[29480] + MEM[30025];
assign MEM[40098] = MEM[29531] + MEM[29688];
assign MEM[40099] = MEM[29553] + MEM[29874];
assign MEM[40100] = MEM[29639] + MEM[29999];
assign MEM[40101] = MEM[29688] + MEM[30251];
assign MEM[40102] = MEM[29694] + MEM[29956];
assign MEM[40103] = MEM[29704] + MEM[29765];
assign MEM[40104] = MEM[29704] + MEM[30101];
assign MEM[40105] = MEM[29708] + MEM[29791];
assign MEM[40106] = MEM[29713] + MEM[29821];
assign MEM[40107] = MEM[29722] + MEM[29797];
assign MEM[40108] = MEM[29723] + MEM[29730];
assign MEM[40109] = MEM[29723] + MEM[29788];
assign MEM[40110] = MEM[29730] + MEM[29821];
assign MEM[40111] = MEM[29733] + MEM[29773];
assign MEM[40112] = MEM[29745] + MEM[29873];
assign MEM[40113] = MEM[29750] + MEM[30065];
assign MEM[40114] = MEM[29763] + MEM[29895];
assign MEM[40115] = MEM[29764] + MEM[29797];
assign MEM[40116] = MEM[29764] + MEM[29841];
assign MEM[40117] = MEM[29765] + MEM[29924];
assign MEM[40118] = MEM[29780] + MEM[29913];
assign MEM[40119] = MEM[29784] + MEM[29829];
assign MEM[40120] = MEM[29786] + MEM[30043];
assign MEM[40121] = MEM[29786] + MEM[30206];
assign MEM[40122] = MEM[29791] + MEM[30294];
assign MEM[40123] = MEM[29793] + MEM[29794];
assign MEM[40124] = MEM[29794] + MEM[30531];
assign MEM[40125] = MEM[29801] + MEM[30120];
assign MEM[40126] = MEM[29811] + MEM[30165];
assign MEM[40127] = MEM[29847] + MEM[29850];
assign MEM[40128] = MEM[29850] + MEM[29888];
assign MEM[40129] = MEM[29857] + MEM[29990];
assign MEM[40130] = MEM[29857] + MEM[30169];
assign MEM[40131] = MEM[29868] + MEM[30075];
assign MEM[40132] = MEM[29868] + MEM[30159];
assign MEM[40133] = MEM[29873] + MEM[29924];
assign MEM[40134] = MEM[29874] + MEM[29999];
assign MEM[40135] = MEM[29885] + MEM[29930];
assign MEM[40136] = MEM[29886] + MEM[29935];
assign MEM[40137] = MEM[29886] + MEM[30277];
assign MEM[40138] = MEM[29888] + MEM[29932];
assign MEM[40139] = MEM[29895] + MEM[30085];
assign MEM[40140] = MEM[29913] + MEM[30664];
assign MEM[40141] = MEM[29914] + MEM[29990];
assign MEM[40142] = MEM[29914] + MEM[30121];
assign MEM[40143] = MEM[29927] + MEM[29950];
assign MEM[40144] = MEM[29927] + MEM[29991];
assign MEM[40145] = MEM[29930] + MEM[30271];
assign MEM[40146] = MEM[29935] + MEM[30457];
assign MEM[40147] = MEM[29938] + MEM[30074];
assign MEM[40148] = MEM[29938] + MEM[30099];
assign MEM[40149] = MEM[29950] + MEM[30074];
assign MEM[40150] = MEM[29956] + MEM[30085];
assign MEM[40151] = MEM[29982] + MEM[30137];
assign MEM[40152] = MEM[29991] + MEM[30121];
assign MEM[40153] = MEM[29993] + MEM[30049];
assign MEM[40154] = MEM[29993] + MEM[30351];
assign MEM[40155] = MEM[30019] + MEM[30322];
assign MEM[40156] = MEM[30022] + MEM[30115];
assign MEM[40157] = MEM[30022] + MEM[30553];
assign MEM[40158] = MEM[30025] + MEM[30075];
assign MEM[40159] = MEM[30027] + MEM[30249];
assign MEM[40160] = MEM[30027] + MEM[30332];
assign MEM[40161] = MEM[30041] + MEM[30115];
assign MEM[40162] = MEM[30041] + MEM[30220];
assign MEM[40163] = MEM[30043] + MEM[30045];
assign MEM[40164] = MEM[30045] + MEM[30290];
assign MEM[40165] = MEM[30046] + MEM[30250];
assign MEM[40166] = MEM[30046] + MEM[30688];
assign MEM[40167] = MEM[30049] + MEM[30263];
assign MEM[40168] = MEM[30050] + MEM[30299];
assign MEM[40169] = MEM[30050] + MEM[30317];
assign MEM[40170] = MEM[30061] + MEM[30258];
assign MEM[40171] = MEM[30099] + MEM[30284];
assign MEM[40172] = MEM[30101] + MEM[30286];
assign MEM[40173] = MEM[30109] + MEM[30158];
assign MEM[40174] = MEM[30109] + MEM[30411];
assign MEM[40175] = MEM[30120] + MEM[30249];
assign MEM[40176] = MEM[30126] + MEM[30220];
assign MEM[40177] = MEM[30126] + MEM[30267];
assign MEM[40178] = MEM[30137] + MEM[30284];
assign MEM[40179] = MEM[30158] + MEM[30159];
assign MEM[40180] = MEM[30162] + MEM[30331];
assign MEM[40181] = MEM[30162] + MEM[30387];
assign MEM[40182] = MEM[30165] + MEM[30238];
assign MEM[40183] = MEM[30169] + MEM[30304];
assign MEM[40184] = MEM[30192] + MEM[30223];
assign MEM[40185] = MEM[30192] + MEM[30338];
assign MEM[40186] = MEM[30205] + MEM[30258];
assign MEM[40187] = MEM[30205] + MEM[30515];
assign MEM[40188] = MEM[30206] + MEM[30447];
assign MEM[40189] = MEM[30207] + MEM[30246];
assign MEM[40190] = MEM[30207] + MEM[30259];
assign MEM[40191] = MEM[30210] + MEM[30235];
assign MEM[40192] = MEM[30210] + MEM[30423];
assign MEM[40193] = MEM[30223] + MEM[30246];
assign MEM[40194] = MEM[30235] + MEM[30441];
assign MEM[40195] = MEM[30236] + MEM[30263];
assign MEM[40196] = MEM[30236] + MEM[30475];
assign MEM[40197] = MEM[30238] + MEM[30825];
assign MEM[40198] = MEM[30250] + MEM[30256];
assign MEM[40199] = MEM[30251] + MEM[30420];
assign MEM[40200] = MEM[30256] + MEM[30311];
assign MEM[40201] = MEM[30259] + MEM[30515];
assign MEM[40202] = MEM[30267] + MEM[30360];
assign MEM[40203] = MEM[30270] + MEM[30298];
assign MEM[40204] = MEM[30270] + MEM[30343];
assign MEM[40205] = MEM[30271] + MEM[30470];
assign MEM[40206] = MEM[30277] + MEM[30341];
assign MEM[40207] = MEM[30286] + MEM[30339];
assign MEM[40208] = MEM[30290] + MEM[30671];
assign MEM[40209] = MEM[30294] + MEM[30468];
assign MEM[40210] = MEM[30298] + MEM[30301];
assign MEM[40211] = MEM[30299] + MEM[30416];
assign MEM[40212] = MEM[30301] + MEM[30311];
assign MEM[40213] = MEM[30304] + MEM[30532];
assign MEM[40214] = MEM[30313] + MEM[30343];
assign MEM[40215] = MEM[30313] + MEM[30398];
assign MEM[40216] = MEM[30317] + MEM[30526];
assign MEM[40217] = MEM[30322] + MEM[30494];
assign MEM[40218] = MEM[30331] + MEM[30441];
assign MEM[40219] = MEM[30332] + MEM[30338];
assign MEM[40220] = MEM[30339] + MEM[30413];
assign MEM[40221] = MEM[30341] + MEM[30554];
assign MEM[40222] = MEM[30351] + MEM[30359];
assign MEM[40223] = MEM[30359] + MEM[30585];
assign MEM[40224] = MEM[30360] + MEM[30406];
assign MEM[40225] = MEM[30365] + MEM[30394];
assign MEM[40226] = MEM[30365] + MEM[30575];
assign MEM[40227] = MEM[30376] + MEM[30419];
assign MEM[40228] = MEM[30376] + MEM[30551];
assign MEM[40229] = MEM[30383] + MEM[30574];
assign MEM[40230] = MEM[30383] + MEM[30864];
assign MEM[40231] = MEM[30387] + MEM[30568];
assign MEM[40232] = MEM[30394] + MEM[30878];
assign MEM[40233] = MEM[30398] + MEM[30874];
assign MEM[40234] = MEM[30406] + MEM[30584];
assign MEM[40235] = MEM[30411] + MEM[30467];
assign MEM[40236] = MEM[30413] + MEM[30642];
assign MEM[40237] = MEM[30416] + MEM[30760];
assign MEM[40238] = MEM[30419] + MEM[30657];
assign MEM[40239] = MEM[30420] + MEM[30617];
assign MEM[40240] = MEM[30423] + MEM[30446];
assign MEM[40241] = MEM[30432] + MEM[30467];
assign MEM[40242] = MEM[30432] + MEM[30809];
assign MEM[40243] = MEM[30446] + MEM[30532];
assign MEM[40244] = MEM[30447] + MEM[30648];
assign MEM[40245] = MEM[30457] + MEM[30480];
assign MEM[40246] = MEM[30468] + MEM[30470];
assign MEM[40247] = MEM[30473] + MEM[30483];
assign MEM[40248] = MEM[30473] + MEM[30617];
assign MEM[40249] = MEM[30475] + MEM[30531];
assign MEM[40250] = MEM[30480] + MEM[30635];
assign MEM[40251] = MEM[30482] + MEM[30510];
assign MEM[40252] = MEM[30482] + MEM[30666];
assign MEM[40253] = MEM[30483] + MEM[30494];
assign MEM[40254] = MEM[30485] + MEM[30580];
assign MEM[40255] = MEM[30485] + MEM[30729];
assign MEM[40256] = MEM[30499] + MEM[30648];
assign MEM[40257] = MEM[30499] + MEM[30665];
assign MEM[40258] = MEM[30510] + MEM[30526];
assign MEM[40259] = MEM[30534] + MEM[30667];
assign MEM[40260] = MEM[30534] + MEM[30708];
assign MEM[40261] = MEM[30551] + MEM[30601];
assign MEM[40262] = MEM[30553] + MEM[30732];
assign MEM[40263] = MEM[30554] + MEM[31009];
assign MEM[40264] = MEM[30556] + MEM[30568];
assign MEM[40265] = MEM[30556] + MEM[30715];
assign MEM[40266] = MEM[30565] + MEM[30773];
assign MEM[40267] = MEM[30565] + MEM[30810];
assign MEM[40268] = MEM[30574] + MEM[30584];
assign MEM[40269] = MEM[30575] + MEM[30635];
assign MEM[40270] = MEM[30580] + MEM[30665];
assign MEM[40271] = MEM[30585] + MEM[30595];
assign MEM[40272] = MEM[30586] + MEM[30640];
assign MEM[40273] = MEM[30586] + MEM[30770];
assign MEM[40274] = MEM[30595] + MEM[30613];
assign MEM[40275] = MEM[30601] + MEM[30791];
assign MEM[40276] = MEM[30606] + MEM[30661];
assign MEM[40277] = MEM[30606] + MEM[30732];
assign MEM[40278] = MEM[30611] + MEM[30657];
assign MEM[40279] = MEM[30611] + MEM[30712];
assign MEM[40280] = MEM[30613] + MEM[30696];
assign MEM[40281] = MEM[30625] + MEM[30881];
assign MEM[40282] = MEM[30625] + MEM[30990];
assign MEM[40283] = MEM[30627] + MEM[30667];
assign MEM[40284] = MEM[30627] + MEM[30846];
assign MEM[40285] = MEM[30640] + MEM[30743];
assign MEM[40286] = MEM[30642] + MEM[30773];
assign MEM[40287] = MEM[30661] + MEM[30881];
assign MEM[40288] = MEM[30664] + MEM[30692];
assign MEM[40289] = MEM[30666] + MEM[30692];
assign MEM[40290] = MEM[30671] + MEM[30725];
assign MEM[40291] = MEM[30675] + MEM[30718];
assign MEM[40292] = MEM[30675] + MEM[30866];
assign MEM[40293] = MEM[30686] + MEM[30698];
assign MEM[40294] = MEM[30686] + MEM[30971];
assign MEM[40295] = MEM[30688] + MEM[30838];
assign MEM[40296] = MEM[30696] + MEM[30720];
assign MEM[40297] = MEM[30698] + MEM[30933];
assign MEM[40298] = MEM[30701] + MEM[30797];
assign MEM[40299] = MEM[30701] + MEM[30905];
assign MEM[40300] = MEM[30704] + MEM[30812];
assign MEM[40301] = MEM[30704] + MEM[30850];
assign MEM[40302] = MEM[30708] + MEM[30829];
assign MEM[40303] = MEM[30712] + MEM[30716];
assign MEM[40304] = MEM[30715] + MEM[30729];
assign MEM[40305] = MEM[30716] + MEM[30977];
assign MEM[40306] = MEM[30718] + MEM[30878];
assign MEM[40307] = MEM[30720] + MEM[30902];
assign MEM[40308] = MEM[30725] + MEM[30825];
assign MEM[40309] = MEM[30734] + MEM[30762];
assign MEM[40310] = MEM[30734] + MEM[31001];
assign MEM[40311] = MEM[30743] + MEM[30928];
assign MEM[40312] = MEM[30746] + MEM[30856];
assign MEM[40313] = MEM[30746] + MEM[31029];
assign MEM[40314] = MEM[30760] + MEM[31001];
assign MEM[40315] = MEM[30762] + MEM[30770];
assign MEM[40316] = MEM[30776] + MEM[30927];
assign MEM[40317] = MEM[30776] + MEM[31056];
assign MEM[40318] = MEM[30784] + MEM[31305];
assign MEM[40319] = MEM[30784] + MEM[31369];
assign MEM[40320] = MEM[30787] + MEM[30834];
assign MEM[40321] = MEM[30787] + MEM[31207];
assign MEM[40322] = MEM[30788] + MEM[30818];
assign MEM[40323] = MEM[30788] + MEM[31060];
assign MEM[40324] = MEM[30791] + MEM[31083];
assign MEM[40325] = MEM[30795] + MEM[30826];
assign MEM[40326] = MEM[30795] + MEM[30940];
assign MEM[40327] = MEM[30797] + MEM[30987];
assign MEM[40328] = MEM[30809] + MEM[30810];
assign MEM[40329] = MEM[30812] + MEM[30983];
assign MEM[40330] = MEM[30813] + MEM[30829];
assign MEM[40331] = MEM[30813] + MEM[30951];
assign MEM[40332] = MEM[30818] + MEM[30923];
assign MEM[40333] = MEM[30826] + MEM[30908];
assign MEM[40334] = MEM[30834] + MEM[30887];
assign MEM[40335] = MEM[30838] + MEM[30902];
assign MEM[40336] = MEM[30844] + MEM[30917];
assign MEM[40337] = MEM[30844] + MEM[31009];
assign MEM[40338] = MEM[30846] + MEM[30932];
assign MEM[40339] = MEM[30849] + MEM[30951];
assign MEM[40340] = MEM[30849] + MEM[31006];
assign MEM[40341] = MEM[30850] + MEM[30856];
assign MEM[40342] = MEM[30852] + MEM[30857];
assign MEM[40343] = MEM[30852] + MEM[30900];
assign MEM[40344] = MEM[30857] + MEM[30997];
assign MEM[40345] = MEM[30864] + MEM[30877];
assign MEM[40346] = MEM[30866] + MEM[30959];
assign MEM[40347] = MEM[30874] + MEM[30908];
assign MEM[40348] = MEM[30877] + MEM[30907];
assign MEM[40349] = MEM[30882] + MEM[30932];
assign MEM[40350] = MEM[30882] + MEM[31212];
assign MEM[40351] = MEM[30887] + MEM[30937];
assign MEM[40352] = MEM[30889] + MEM[30966];
assign MEM[40353] = MEM[30889] + MEM[31175];
assign MEM[40354] = MEM[30900] + MEM[30917];
assign MEM[40355] = MEM[30905] + MEM[30927];
assign MEM[40356] = MEM[30907] + MEM[31098];
assign MEM[40357] = MEM[30915] + MEM[30928];
assign MEM[40358] = MEM[30915] + MEM[30952];
assign MEM[40359] = MEM[30923] + MEM[30940];
assign MEM[40360] = MEM[30933] + MEM[30952];
assign MEM[40361] = MEM[30937] + MEM[30958];
assign MEM[40362] = MEM[30939] + MEM[30942];
assign MEM[40363] = MEM[30939] + MEM[31139];
assign MEM[40364] = MEM[30941] + MEM[30977];
assign MEM[40365] = MEM[30941] + MEM[30981];
assign MEM[40366] = MEM[30942] + MEM[31269];
assign MEM[40367] = MEM[30958] + MEM[31023];
assign MEM[40368] = MEM[30959] + MEM[31276];
assign MEM[40369] = MEM[30966] + MEM[30999];
assign MEM[40370] = MEM[30971] + MEM[31089];
assign MEM[40371] = MEM[30981] + MEM[31129];
assign MEM[40372] = MEM[30983] + MEM[30999];
assign MEM[40373] = MEM[30985] + MEM[31084];
assign MEM[40374] = MEM[30985] + MEM[31127];
assign MEM[40375] = MEM[30987] + MEM[31400];
assign MEM[40376] = MEM[30990] + MEM[31131];
assign MEM[40377] = MEM[30991] + MEM[31039];
assign MEM[40378] = MEM[30991] + MEM[31252];
assign MEM[40379] = MEM[30997] + MEM[31061];
assign MEM[40380] = MEM[31006] + MEM[31018];
assign MEM[40381] = MEM[31011] + MEM[31014];
assign MEM[40382] = MEM[31011] + MEM[31284];
assign MEM[40383] = MEM[31014] + MEM[31279];
assign MEM[40384] = MEM[31018] + MEM[31147];
assign MEM[40385] = MEM[31023] + MEM[31357];
assign MEM[40386] = MEM[31029] + MEM[31083];
assign MEM[40387] = MEM[31039] + MEM[31536];
assign MEM[40388] = MEM[31045] + MEM[31174];
assign MEM[40389] = MEM[31045] + MEM[31189];
assign MEM[40390] = MEM[31046] + MEM[31061];
assign MEM[40391] = MEM[31046] + MEM[31164];
assign MEM[40392] = MEM[31048] + MEM[31063];
assign MEM[40393] = MEM[31048] + MEM[31261];
assign MEM[40394] = MEM[31056] + MEM[31153];
assign MEM[40395] = MEM[31060] + MEM[31334];
assign MEM[40396] = MEM[31063] + MEM[31205];
assign MEM[40397] = MEM[31071] + MEM[31235];
assign MEM[40398] = MEM[31071] + MEM[31245];
assign MEM[40399] = MEM[31074] + MEM[31203];
assign MEM[40400] = MEM[31074] + MEM[31235];
assign MEM[40401] = MEM[31078] + MEM[31281];
assign MEM[40402] = MEM[31078] + MEM[31383];
assign MEM[40403] = MEM[31084] + MEM[31207];
assign MEM[40404] = MEM[31089] + MEM[31144];
assign MEM[40405] = MEM[31095] + MEM[31107];
assign MEM[40406] = MEM[31095] + MEM[31265];
assign MEM[40407] = MEM[31098] + MEM[31409];
assign MEM[40408] = MEM[31106] + MEM[31151];
assign MEM[40409] = MEM[31106] + MEM[31341];
assign MEM[40410] = MEM[31107] + MEM[31164];
assign MEM[40411] = MEM[31112] + MEM[31205];
assign MEM[40412] = MEM[31112] + MEM[31409];
assign MEM[40413] = MEM[31120] + MEM[31223];
assign MEM[40414] = MEM[31120] + MEM[31248];
assign MEM[40415] = MEM[31127] + MEM[31139];
assign MEM[40416] = MEM[31129] + MEM[31444];
assign MEM[40417] = MEM[31131] + MEM[31373];
assign MEM[40418] = MEM[31144] + MEM[31183];
assign MEM[40419] = MEM[31147] + MEM[31151];
assign MEM[40420] = MEM[31153] + MEM[31278];
assign MEM[40421] = MEM[31173] + MEM[31183];
assign MEM[40422] = MEM[31173] + MEM[31213];
assign MEM[40423] = MEM[31174] + MEM[31494];
assign MEM[40424] = MEM[31175] + MEM[31344];
assign MEM[40425] = MEM[31176] + MEM[31237];
assign MEM[40426] = MEM[31176] + MEM[31285];
assign MEM[40427] = MEM[31188] + MEM[31189];
assign MEM[40428] = MEM[31188] + MEM[31331];
assign MEM[40429] = MEM[31203] + MEM[31248];
assign MEM[40430] = MEM[31209] + MEM[31213];
assign MEM[40431] = MEM[31209] + MEM[31261];
assign MEM[40432] = MEM[31212] + MEM[31329];
assign MEM[40433] = MEM[31214] + MEM[31221];
assign MEM[40434] = MEM[31214] + MEM[31291];
assign MEM[40435] = MEM[31221] + MEM[31246];
assign MEM[40436] = MEM[31223] + MEM[31447];
assign MEM[40437] = MEM[31225] + MEM[31252];
assign MEM[40438] = MEM[31225] + MEM[31379];
assign MEM[40439] = MEM[31228] + MEM[31303];
assign MEM[40440] = MEM[31228] + MEM[31375];
assign MEM[40441] = MEM[31237] + MEM[31281];
assign MEM[40442] = MEM[31238] + MEM[31244];
assign MEM[40443] = MEM[31238] + MEM[31327];
assign MEM[40444] = MEM[31244] + MEM[31269];
assign MEM[40445] = MEM[31245] + MEM[31429];
assign MEM[40446] = MEM[31246] + MEM[31341];
assign MEM[40447] = MEM[31265] + MEM[31374];
assign MEM[40448] = MEM[31270] + MEM[31324];
assign MEM[40449] = MEM[31270] + MEM[31600];
assign MEM[40450] = MEM[31276] + MEM[31279];
assign MEM[40451] = MEM[31277] + MEM[31293];
assign MEM[40452] = MEM[31277] + MEM[31483];
assign MEM[40453] = MEM[31278] + MEM[31299];
assign MEM[40454] = MEM[31283] + MEM[31311];
assign MEM[40455] = MEM[31283] + MEM[31379];
assign MEM[40456] = MEM[31284] + MEM[31299];
assign MEM[40457] = MEM[31285] + MEM[31305];
assign MEM[40458] = MEM[31288] + MEM[31291];
assign MEM[40459] = MEM[31288] + MEM[31453];
assign MEM[40460] = MEM[31293] + MEM[31357];
assign MEM[40461] = MEM[31303] + MEM[31586];
assign MEM[40462] = MEM[31311] + MEM[31403];
assign MEM[40463] = MEM[31324] + MEM[31334];
assign MEM[40464] = MEM[31327] + MEM[31441];
assign MEM[40465] = MEM[31329] + MEM[31407];
assign MEM[40466] = MEM[31331] + MEM[31452];
assign MEM[40467] = MEM[31335] + MEM[31362];
assign MEM[40468] = MEM[31335] + MEM[31374];
assign MEM[40469] = MEM[31343] + MEM[31362];
assign MEM[40470] = MEM[31343] + MEM[31469];
assign MEM[40471] = MEM[31344] + MEM[31407];
assign MEM[40472] = MEM[31345] + MEM[31460];
assign MEM[40473] = MEM[31345] + MEM[31586];
assign MEM[40474] = MEM[31348] + MEM[31416];
assign MEM[40475] = MEM[31348] + MEM[31749];
assign MEM[40476] = MEM[31350] + MEM[31378];
assign MEM[40477] = MEM[31350] + MEM[31420];
assign MEM[40478] = MEM[31359] + MEM[31452];
assign MEM[40479] = MEM[31359] + MEM[31484];
assign MEM[40480] = MEM[31369] + MEM[31497];
assign MEM[40481] = MEM[31373] + MEM[31416];
assign MEM[40482] = MEM[31375] + MEM[31651];
assign MEM[40483] = MEM[31378] + MEM[31504];
assign MEM[40484] = MEM[31383] + MEM[31417];
assign MEM[40485] = MEM[31385] + MEM[31417];
assign MEM[40486] = MEM[31385] + MEM[31676];
assign MEM[40487] = MEM[31389] + MEM[31394];
assign MEM[40488] = MEM[31389] + MEM[31672];
assign MEM[40489] = MEM[31394] + MEM[31441];
assign MEM[40490] = MEM[31400] + MEM[31435];
assign MEM[40491] = MEM[31403] + MEM[31457];
assign MEM[40492] = MEM[31404] + MEM[31440];
assign MEM[40493] = MEM[31404] + MEM[31499];
assign MEM[40494] = MEM[31412] + MEM[31413];
assign MEM[40495] = MEM[31412] + MEM[31692];
assign MEM[40496] = MEM[31413] + MEM[31471];
assign MEM[40497] = MEM[31418] + MEM[31431];
assign MEM[40498] = MEM[31418] + MEM[31437];
assign MEM[40499] = MEM[31420] + MEM[31500];
assign MEM[40500] = MEM[31429] + MEM[31453];
assign MEM[40501] = MEM[31431] + MEM[31435];
assign MEM[40502] = MEM[31437] + MEM[31478];
assign MEM[40503] = MEM[31440] + MEM[31457];
assign MEM[40504] = MEM[31444] + MEM[31756];
assign MEM[40505] = MEM[31447] + MEM[31459];
assign MEM[40506] = MEM[31456] + MEM[31520];
assign MEM[40507] = MEM[31456] + MEM[31537];
assign MEM[40508] = MEM[31459] + MEM[31545];
assign MEM[40509] = MEM[31460] + MEM[31546];
assign MEM[40510] = MEM[31468] + MEM[31479];
assign MEM[40511] = MEM[31468] + MEM[31590];
assign MEM[40512] = MEM[31469] + MEM[31685];
assign MEM[40513] = MEM[31471] + MEM[31584];
assign MEM[40514] = MEM[31478] + MEM[31549];
assign MEM[40515] = MEM[31479] + MEM[31490];
assign MEM[40516] = MEM[31483] + MEM[31667];
assign MEM[40517] = MEM[31484] + MEM[31594];
assign MEM[40518] = MEM[31490] + MEM[31584];
assign MEM[40519] = MEM[31494] + MEM[31673];
assign MEM[40520] = MEM[31497] + MEM[31596];
assign MEM[40521] = MEM[31499] + MEM[31568];
assign MEM[40522] = MEM[31500] + MEM[31554];
assign MEM[40523] = MEM[31504] + MEM[31525];
assign MEM[40524] = MEM[31511] + MEM[31607];
assign MEM[40525] = MEM[31511] + MEM[31617];
assign MEM[40526] = MEM[31520] + MEM[31550];
assign MEM[40527] = MEM[31524] + MEM[31617];
assign MEM[40528] = MEM[31524] + MEM[31756];
assign MEM[40529] = MEM[31525] + MEM[31616];
assign MEM[40530] = MEM[31529] + MEM[31537];
assign MEM[40531] = MEM[31529] + MEM[31538];
assign MEM[40532] = MEM[31536] + MEM[31544];
assign MEM[40533] = MEM[31538] + MEM[31753];
assign MEM[40534] = MEM[31544] + MEM[31758];
assign MEM[40535] = MEM[31545] + MEM[31633];
assign MEM[40536] = MEM[31546] + MEM[31572];
assign MEM[40537] = MEM[31549] + MEM[31731];
assign MEM[40538] = MEM[31550] + MEM[31565];
assign MEM[40539] = MEM[31551] + MEM[31596];
assign MEM[40540] = MEM[31551] + MEM[31599];
assign MEM[40541] = MEM[31552] + MEM[31703];
assign MEM[40542] = MEM[31552] + MEM[31725];
assign MEM[40543] = MEM[31554] + MEM[31662];
assign MEM[40544] = MEM[31562] + MEM[31572];
assign MEM[40545] = MEM[31562] + MEM[31746];
assign MEM[40546] = MEM[31563] + MEM[31593];
assign MEM[40547] = MEM[31563] + MEM[31669];
assign MEM[40548] = MEM[31565] + MEM[31602];
assign MEM[40549] = MEM[31568] + MEM[31634];
assign MEM[40550] = MEM[31590] + MEM[31602];
assign MEM[40551] = MEM[31593] + MEM[31597];
assign MEM[40552] = MEM[31594] + MEM[31722];
assign MEM[40553] = MEM[31597] + MEM[31613];
assign MEM[40554] = MEM[31599] + MEM[31650];
assign MEM[40555] = MEM[31600] + MEM[31796];
assign MEM[40556] = MEM[31607] + MEM[31760];
assign MEM[40557] = MEM[31610] + MEM[31672];
assign MEM[40558] = MEM[31610] + MEM[31732];
assign MEM[40559] = MEM[31613] + MEM[31614];
assign MEM[40560] = MEM[31614] + MEM[31619];
assign MEM[40561] = MEM[31616] + MEM[31749];
assign MEM[40562] = MEM[31619] + MEM[31633];
assign MEM[40563] = MEM[31620] + MEM[31637];
assign MEM[40564] = MEM[31620] + MEM[31641];
assign MEM[40565] = MEM[31627] + MEM[31634];
assign MEM[40566] = MEM[31627] + MEM[31827];
assign MEM[40567] = MEM[31637] + MEM[31663];
assign MEM[40568] = MEM[31641] + MEM[31951];
assign MEM[40569] = MEM[31644] + MEM[31645];
assign MEM[40570] = MEM[31644] + MEM[31667];
assign MEM[40571] = MEM[31645] + MEM[31965];
assign MEM[40572] = MEM[31650] + MEM[31664];
assign MEM[40573] = MEM[31651] + MEM[32027];
assign MEM[40574] = MEM[31655] + MEM[31740];
assign MEM[40575] = MEM[31655] + MEM[31770];
assign MEM[40576] = MEM[31657] + MEM[31663];
assign MEM[40577] = MEM[31657] + MEM[31673];
assign MEM[40578] = MEM[31662] + MEM[31664];
assign MEM[40579] = MEM[31666] + MEM[31704];
assign MEM[40580] = MEM[31666] + MEM[31829];
assign MEM[40581] = MEM[31669] + MEM[31789];
assign MEM[40582] = MEM[31676] + MEM[31703];
assign MEM[40583] = MEM[31683] + MEM[31701];
assign MEM[40584] = MEM[31683] + MEM[31738];
assign MEM[40585] = MEM[31685] + MEM[31787];
assign MEM[40586] = MEM[31692] + MEM[31783];
assign MEM[40587] = MEM[31701] + MEM[31714];
assign MEM[40588] = MEM[31704] + MEM[32251];
assign MEM[40589] = MEM[31706] + MEM[31787];
assign MEM[40590] = MEM[31706] + MEM[32107];
assign MEM[40591] = MEM[31713] + MEM[31783];
assign MEM[40592] = MEM[31713] + MEM[31939];
assign MEM[40593] = MEM[31714] + MEM[31852];
assign MEM[40594] = MEM[31721] + MEM[31732];
assign MEM[40595] = MEM[31721] + MEM[31746];
assign MEM[40596] = MEM[31722] + MEM[31843];
assign MEM[40597] = MEM[31723] + MEM[31725];
assign MEM[40598] = MEM[31723] + MEM[31784];
assign MEM[40599] = MEM[31731] + MEM[31736];
assign MEM[40600] = MEM[31736] + MEM[31784];
assign MEM[40601] = MEM[31738] + MEM[31798];
assign MEM[40602] = MEM[31740] + MEM[31791];
assign MEM[40603] = MEM[31747] + MEM[31774];
assign MEM[40604] = MEM[31747] + MEM[31812];
assign MEM[40605] = MEM[31752] + MEM[31761];
assign MEM[40606] = MEM[31752] + MEM[31815];
assign MEM[40607] = MEM[31753] + MEM[31760];
assign MEM[40608] = MEM[31758] + MEM[31930];
assign MEM[40609] = MEM[31761] + MEM[31999];
assign MEM[40610] = MEM[31770] + MEM[31819];
assign MEM[40611] = MEM[31774] + MEM[32007];
assign MEM[40612] = MEM[31775] + MEM[31788];
assign MEM[40613] = MEM[31775] + MEM[31789];
assign MEM[40614] = MEM[31778] + MEM[31782];
assign MEM[40615] = MEM[31778] + MEM[32070];
assign MEM[40616] = MEM[31782] + MEM[31826];
assign MEM[40617] = MEM[31788] + MEM[31794];
assign MEM[40618] = MEM[31791] + MEM[31815];
assign MEM[40619] = MEM[31793] + MEM[31837];
assign MEM[40620] = MEM[31793] + MEM[31861];
assign MEM[40621] = MEM[31794] + MEM[31801];
assign MEM[40622] = MEM[31796] + MEM[32131];
assign MEM[40623] = MEM[31798] + MEM[31812];
assign MEM[40624] = MEM[31801] + MEM[31997];
assign MEM[40625] = MEM[31802] + MEM[31807];
assign MEM[40626] = MEM[31802] + MEM[31811];
assign MEM[40627] = MEM[31807] + MEM[31814];
assign MEM[40628] = MEM[31810] + MEM[31950];
assign MEM[40629] = MEM[31810] + MEM[31970];
assign MEM[40630] = MEM[31811] + MEM[31905];
assign MEM[40631] = MEM[31814] + MEM[31971];
assign MEM[40632] = MEM[31816] + MEM[31887];
assign MEM[40633] = MEM[31816] + MEM[32138];
assign MEM[40634] = MEM[31819] + MEM[31876];
assign MEM[40635] = MEM[31820] + MEM[31822];
assign MEM[40636] = MEM[31820] + MEM[31843];
assign MEM[40637] = MEM[31822] + MEM[31995];
assign MEM[40638] = MEM[31826] + MEM[31883];
assign MEM[40639] = MEM[31827] + MEM[31935];
assign MEM[40640] = MEM[31829] + MEM[31889];
assign MEM[40641] = MEM[31831] + MEM[31883];
assign MEM[40642] = MEM[31831] + MEM[32003];
assign MEM[40643] = MEM[31834] + MEM[31863];
assign MEM[40644] = MEM[31834] + MEM[32014];
assign MEM[40645] = MEM[31837] + MEM[31885];
assign MEM[40646] = MEM[31841] + MEM[31866];
assign MEM[40647] = MEM[31841] + MEM[31995];
assign MEM[40648] = MEM[31852] + MEM[31896];
assign MEM[40649] = MEM[31861] + MEM[31944];
assign MEM[40650] = MEM[31862] + MEM[31882];
assign MEM[40651] = MEM[31862] + MEM[32007];
assign MEM[40652] = MEM[31863] + MEM[31887];
assign MEM[40653] = MEM[31866] + MEM[31897];
assign MEM[40654] = MEM[31876] + MEM[32132];
assign MEM[40655] = MEM[31881] + MEM[32040];
assign MEM[40656] = MEM[31881] + MEM[32075];
assign MEM[40657] = MEM[31882] + MEM[31965];
assign MEM[40658] = MEM[31885] + MEM[32044];
assign MEM[40659] = MEM[31889] + MEM[32014];
assign MEM[40660] = MEM[31890] + MEM[31910];
assign MEM[40661] = MEM[31890] + MEM[31958];
assign MEM[40662] = MEM[31896] + MEM[32003];
assign MEM[40663] = MEM[31897] + MEM[31980];
assign MEM[40664] = MEM[31900] + MEM[31920];
assign MEM[40665] = MEM[31900] + MEM[32067];
assign MEM[40666] = MEM[31905] + MEM[31939];
assign MEM[40667] = MEM[31906] + MEM[31909];
assign MEM[40668] = MEM[31906] + MEM[31930];
assign MEM[40669] = MEM[31909] + MEM[32232];
assign MEM[40670] = MEM[31910] + MEM[32054];
assign MEM[40671] = MEM[31920] + MEM[32040];
assign MEM[40672] = MEM[31927] + MEM[31986];
assign MEM[40673] = MEM[31927] + MEM[32021];
assign MEM[40674] = MEM[31934] + MEM[31944];
assign MEM[40675] = MEM[31934] + MEM[31957];
assign MEM[40676] = MEM[31935] + MEM[32059];
assign MEM[40677] = MEM[31942] + MEM[32073];
assign MEM[40678] = MEM[31942] + MEM[32096];
assign MEM[40679] = MEM[31950] + MEM[31957];
assign MEM[40680] = MEM[31951] + MEM[32018];
assign MEM[40681] = MEM[31958] + MEM[32043];
assign MEM[40682] = MEM[31959] + MEM[32085];
assign MEM[40683] = MEM[31959] + MEM[32101];
assign MEM[40684] = MEM[31970] + MEM[31999];
assign MEM[40685] = MEM[31971] + MEM[31986];
assign MEM[40686] = MEM[31972] + MEM[32072];
assign MEM[40687] = MEM[31972] + MEM[32157];
assign MEM[40688] = MEM[31976] + MEM[31991];
assign MEM[40689] = MEM[31976] + MEM[32109];
assign MEM[40690] = MEM[31980] + MEM[32066];
assign MEM[40691] = MEM[31985] + MEM[31998];
assign MEM[40692] = MEM[31985] + MEM[32049];
assign MEM[40693] = MEM[31991] + MEM[31998];
assign MEM[40694] = MEM[31997] + MEM[32043];
assign MEM[40695] = MEM[32001] + MEM[32087];
assign MEM[40696] = MEM[32001] + MEM[32269];
assign MEM[40697] = MEM[32016] + MEM[32049];
assign MEM[40698] = MEM[32016] + MEM[32185];
assign MEM[40699] = MEM[32018] + MEM[32114];
assign MEM[40700] = MEM[32021] + MEM[32078];
assign MEM[40701] = MEM[32027] + MEM[32123];
assign MEM[40702] = MEM[32034] + MEM[32080];
assign MEM[40703] = MEM[32034] + MEM[32221];
assign MEM[40704] = MEM[32044] + MEM[32238];
assign MEM[40705] = MEM[32054] + MEM[32283];
assign MEM[40706] = MEM[32058] + MEM[32188];
assign MEM[40707] = MEM[32058] + MEM[32247];
assign MEM[40708] = MEM[32059] + MEM[32105];
assign MEM[40709] = MEM[32062] + MEM[32131];
assign MEM[40710] = MEM[32062] + MEM[32304];
assign MEM[40711] = MEM[32066] + MEM[32336];
assign MEM[40712] = MEM[32067] + MEM[32088];
assign MEM[40713] = MEM[32070] + MEM[32200];
assign MEM[40714] = MEM[32072] + MEM[32115];
assign MEM[40715] = MEM[32073] + MEM[32237];
assign MEM[40716] = MEM[32075] + MEM[32087];
assign MEM[40717] = MEM[32078] + MEM[32101];
assign MEM[40718] = MEM[32079] + MEM[32092];
assign MEM[40719] = MEM[32079] + MEM[32176];
assign MEM[40720] = MEM[32080] + MEM[32090];
assign MEM[40721] = MEM[32085] + MEM[32089];
assign MEM[40722] = MEM[32088] + MEM[32190];
assign MEM[40723] = MEM[32089] + MEM[32142];
assign MEM[40724] = MEM[32090] + MEM[32149];
assign MEM[40725] = MEM[32092] + MEM[32381];
assign MEM[40726] = MEM[32096] + MEM[32190];
assign MEM[40727] = MEM[32105] + MEM[32200];
assign MEM[40728] = MEM[32107] + MEM[32248];
assign MEM[40729] = MEM[32109] + MEM[32250];
assign MEM[40730] = MEM[32114] + MEM[32132];
assign MEM[40731] = MEM[32115] + MEM[32180];
assign MEM[40732] = MEM[32123] + MEM[32236];
assign MEM[40733] = MEM[32135] + MEM[32139];
assign MEM[40734] = MEM[32135] + MEM[32157];
assign MEM[40735] = MEM[32136] + MEM[32140];
assign MEM[40736] = MEM[32136] + MEM[32343];
assign MEM[40737] = MEM[32138] + MEM[32388];
assign MEM[40738] = MEM[32139] + MEM[32176];
assign MEM[40739] = MEM[32140] + MEM[32166];
assign MEM[40740] = MEM[32142] + MEM[32186];
assign MEM[40741] = MEM[32149] + MEM[32171];
assign MEM[40742] = MEM[32154] + MEM[32166];
assign MEM[40743] = MEM[32154] + MEM[32244];
assign MEM[40744] = MEM[32158] + MEM[32298];
assign MEM[40745] = MEM[32158] + MEM[32343];
assign MEM[40746] = MEM[32171] + MEM[32204];
assign MEM[40747] = MEM[32180] + MEM[32191];
assign MEM[40748] = MEM[32182] + MEM[32400];
assign MEM[40749] = MEM[32182] + MEM[32465];
assign MEM[40750] = MEM[32185] + MEM[32395];
assign MEM[40751] = MEM[32186] + MEM[32252];
assign MEM[40752] = MEM[32188] + MEM[32196];
assign MEM[40753] = MEM[32191] + MEM[32254];
assign MEM[40754] = MEM[32192] + MEM[32198];
assign MEM[40755] = MEM[32192] + MEM[32367];
assign MEM[40756] = MEM[32196] + MEM[32238];
assign MEM[40757] = MEM[32197] + MEM[32214];
assign MEM[40758] = MEM[32197] + MEM[32386];
assign MEM[40759] = MEM[32198] + MEM[32266];
assign MEM[40760] = MEM[32204] + MEM[32242];
assign MEM[40761] = MEM[32208] + MEM[32271];
assign MEM[40762] = MEM[32208] + MEM[32337];
assign MEM[40763] = MEM[32212] + MEM[32308];
assign MEM[40764] = MEM[32212] + MEM[32350];
assign MEM[40765] = MEM[32214] + MEM[32259];
assign MEM[40766] = MEM[32220] + MEM[32250];
assign MEM[40767] = MEM[32220] + MEM[32505];
assign MEM[40768] = MEM[32221] + MEM[32273];
assign MEM[40769] = MEM[32232] + MEM[32311];
assign MEM[40770] = MEM[32236] + MEM[32359];
assign MEM[40771] = MEM[32237] + MEM[32307];
assign MEM[40772] = MEM[32241] + MEM[32251];
assign MEM[40773] = MEM[32241] + MEM[32310];
assign MEM[40774] = MEM[32242] + MEM[32304];
assign MEM[40775] = MEM[32243] + MEM[32261];
assign MEM[40776] = MEM[32243] + MEM[32347];
assign MEM[40777] = MEM[32244] + MEM[32273];
assign MEM[40778] = MEM[32247] + MEM[32259];
assign MEM[40779] = MEM[32248] + MEM[32363];
assign MEM[40780] = MEM[32252] + MEM[32335];
assign MEM[40781] = MEM[32254] + MEM[32282];
assign MEM[40782] = MEM[32261] + MEM[32269];
assign MEM[40783] = MEM[32266] + MEM[32271];
assign MEM[40784] = MEM[32282] + MEM[32306];
assign MEM[40785] = MEM[32283] + MEM[32324];
assign MEM[40786] = MEM[32297] + MEM[32458];
assign MEM[40787] = MEM[32297] + MEM[32533];
assign MEM[40788] = MEM[32298] + MEM[32344];
assign MEM[40789] = MEM[32302] + MEM[32311];
assign MEM[40790] = MEM[32302] + MEM[32733];
assign MEM[40791] = MEM[32306] + MEM[32467];
assign MEM[40792] = MEM[32307] + MEM[32313];
assign MEM[40793] = MEM[32308] + MEM[32338];
assign MEM[40794] = MEM[32309] + MEM[32402];
assign MEM[40795] = MEM[32309] + MEM[32445];
assign MEM[40796] = MEM[32310] + MEM[32335];
assign MEM[40797] = MEM[32313] + MEM[32424];
assign MEM[40798] = MEM[32315] + MEM[32345];
assign MEM[40799] = MEM[32315] + MEM[32497];
assign MEM[40800] = MEM[32317] + MEM[32321];
assign MEM[40801] = MEM[32317] + MEM[32347];
assign MEM[40802] = MEM[32321] + MEM[32506];
assign MEM[40803] = MEM[32324] + MEM[32372];
assign MEM[40804] = MEM[32327] + MEM[32340];
assign MEM[40805] = MEM[32327] + MEM[32397];
assign MEM[40806] = MEM[32336] + MEM[32404];
assign MEM[40807] = MEM[32337] + MEM[32434];
assign MEM[40808] = MEM[32338] + MEM[32392];
assign MEM[40809] = MEM[32340] + MEM[32367];
assign MEM[40810] = MEM[32344] + MEM[32359];
assign MEM[40811] = MEM[32345] + MEM[32612];
assign MEM[40812] = MEM[32350] + MEM[32469];
assign MEM[40813] = MEM[32353] + MEM[32402];
assign MEM[40814] = MEM[32353] + MEM[32405];
assign MEM[40815] = MEM[32355] + MEM[32388];
assign MEM[40816] = MEM[32355] + MEM[32658];
assign MEM[40817] = MEM[32357] + MEM[32375];
assign MEM[40818] = MEM[32357] + MEM[32404];
assign MEM[40819] = MEM[32363] + MEM[32371];
assign MEM[40820] = MEM[32369] + MEM[32464];
assign MEM[40821] = MEM[32369] + MEM[32500];
assign MEM[40822] = MEM[32370] + MEM[32385];
assign MEM[40823] = MEM[32370] + MEM[32400];
assign MEM[40824] = MEM[32371] + MEM[32432];
assign MEM[40825] = MEM[32372] + MEM[32486];
assign MEM[40826] = MEM[32375] + MEM[32453];
assign MEM[40827] = MEM[32379] + MEM[32381];
assign MEM[40828] = MEM[32379] + MEM[32535];
assign MEM[40829] = MEM[32383] + MEM[32410];
assign MEM[40830] = MEM[32383] + MEM[32425];
assign MEM[40831] = MEM[32385] + MEM[32521];
assign MEM[40832] = MEM[32386] + MEM[32398];
assign MEM[40833] = MEM[32392] + MEM[32427];
assign MEM[40834] = MEM[32395] + MEM[32486];
assign MEM[40835] = MEM[32397] + MEM[32450];
assign MEM[40836] = MEM[32398] + MEM[32415];
assign MEM[40837] = MEM[32405] + MEM[32408];
assign MEM[40838] = MEM[32408] + MEM[32473];
assign MEM[40839] = MEM[32410] + MEM[32566];
assign MEM[40840] = MEM[32415] + MEM[32416];
assign MEM[40841] = MEM[32416] + MEM[32614];
assign MEM[40842] = MEM[32419] + MEM[32524];
assign MEM[40843] = MEM[32419] + MEM[32545];
assign MEM[40844] = MEM[32422] + MEM[32443];
assign MEM[40845] = MEM[32422] + MEM[32508];
assign MEM[40846] = MEM[32424] + MEM[32651];
assign MEM[40847] = MEM[32425] + MEM[32474];
assign MEM[40848] = MEM[32427] + MEM[32469];
assign MEM[40849] = MEM[32432] + MEM[32493];
assign MEM[40850] = MEM[32434] + MEM[32454];
assign MEM[40851] = MEM[32443] + MEM[32597];
assign MEM[40852] = MEM[32445] + MEM[32450];
assign MEM[40853] = MEM[32446] + MEM[32517];
assign MEM[40854] = MEM[32446] + MEM[32528];
assign MEM[40855] = MEM[32453] + MEM[32628];
assign MEM[40856] = MEM[32454] + MEM[32479];
assign MEM[40857] = MEM[32458] + MEM[32465];
assign MEM[40858] = MEM[32461] + MEM[32494];
assign MEM[40859] = MEM[32461] + MEM[32583];
assign MEM[40860] = MEM[32464] + MEM[32487];
assign MEM[40861] = MEM[32467] + MEM[32487];
assign MEM[40862] = MEM[32473] + MEM[32566];
assign MEM[40863] = MEM[32474] + MEM[32494];
assign MEM[40864] = MEM[32479] + MEM[32519];
assign MEM[40865] = MEM[32480] + MEM[32501];
assign MEM[40866] = MEM[32480] + MEM[32511];
assign MEM[40867] = MEM[32483] + MEM[32496];
assign MEM[40868] = MEM[32483] + MEM[32700];
assign MEM[40869] = MEM[32490] + MEM[32508];
assign MEM[40870] = MEM[32490] + MEM[32580];
assign MEM[40871] = MEM[32493] + MEM[32516];
assign MEM[40872] = MEM[32495] + MEM[32511];
assign MEM[40873] = MEM[32495] + MEM[32586];
assign MEM[40874] = MEM[32496] + MEM[32516];
assign MEM[40875] = MEM[32497] + MEM[32556];
assign MEM[40876] = MEM[32500] + MEM[32547];
assign MEM[40877] = MEM[32501] + MEM[32540];
assign MEM[40878] = MEM[32505] + MEM[32519];
assign MEM[40879] = MEM[32506] + MEM[32536];
assign MEM[40880] = MEM[32514] + MEM[32545];
assign MEM[40881] = MEM[32514] + MEM[32621];
assign MEM[40882] = MEM[32517] + MEM[32571];
assign MEM[40883] = MEM[32521] + MEM[32534];
assign MEM[40884] = MEM[32523] + MEM[32614];
assign MEM[40885] = MEM[32523] + MEM[32681];
assign MEM[40886] = MEM[32524] + MEM[32535];
assign MEM[40887] = MEM[32527] + MEM[32542];
assign MEM[40888] = MEM[32527] + MEM[32650];
assign MEM[40889] = MEM[32528] + MEM[32548];
assign MEM[40890] = MEM[32531] + MEM[32557];
assign MEM[40891] = MEM[32531] + MEM[32660];
assign MEM[40892] = MEM[32533] + MEM[32607];
assign MEM[40893] = MEM[32534] + MEM[32552];
assign MEM[40894] = MEM[32536] + MEM[32579];
assign MEM[40895] = MEM[32540] + MEM[32558];
assign MEM[40896] = MEM[32542] + MEM[32579];
assign MEM[40897] = MEM[32547] + MEM[32572];
assign MEM[40898] = MEM[32548] + MEM[32602];
assign MEM[40899] = MEM[32552] + MEM[32798];
assign MEM[40900] = MEM[32556] + MEM[32586];
assign MEM[40901] = MEM[32557] + MEM[32564];
assign MEM[40902] = MEM[32558] + MEM[32585];
assign MEM[40903] = MEM[32561] + MEM[32575];
assign MEM[40904] = MEM[32561] + MEM[32613];
assign MEM[40905] = MEM[32564] + MEM[32691];
assign MEM[40906] = MEM[32565] + MEM[32621];
assign MEM[40907] = MEM[32565] + MEM[32954];
assign MEM[40908] = MEM[32570] + MEM[32576];
assign MEM[40909] = MEM[32570] + MEM[32719];
assign MEM[40910] = MEM[32571] + MEM[32667];
assign MEM[40911] = MEM[32572] + MEM[32717];
assign MEM[40912] = MEM[32575] + MEM[32685];
assign MEM[40913] = MEM[32576] + MEM[32666];
assign MEM[40914] = MEM[32577] + MEM[32679];
assign MEM[40915] = MEM[32577] + MEM[32682];
assign MEM[40916] = MEM[32580] + MEM[32646];
assign MEM[40917] = MEM[32583] + MEM[32655];
assign MEM[40918] = MEM[32585] + MEM[32691];
assign MEM[40919] = MEM[32589] + MEM[32593];
assign MEM[40920] = MEM[32589] + MEM[32674];
assign MEM[40921] = MEM[32593] + MEM[32604];
assign MEM[40922] = MEM[32597] + MEM[32738];
assign MEM[40923] = MEM[32602] + MEM[32702];
assign MEM[40924] = MEM[32604] + MEM[32657];
assign MEM[40925] = MEM[32606] + MEM[32613];
assign MEM[40926] = MEM[32606] + MEM[32763];
assign MEM[40927] = MEM[32607] + MEM[32677];
assign MEM[40928] = MEM[32612] + MEM[32658];
assign MEM[40929] = MEM[32615] + MEM[32626];
assign MEM[40930] = MEM[32615] + MEM[32635];
assign MEM[40931] = MEM[32623] + MEM[32662];
assign MEM[40932] = MEM[32623] + MEM[32729];
assign MEM[40933] = MEM[32626] + MEM[32679];
assign MEM[40934] = MEM[32628] + MEM[32635];
assign MEM[40935] = MEM[32646] + MEM[32707];
assign MEM[40936] = MEM[32647] + MEM[32655];
assign MEM[40937] = MEM[32647] + MEM[32668];
assign MEM[40938] = MEM[32649] + MEM[32651];
assign MEM[40939] = MEM[32649] + MEM[32654];
assign MEM[40940] = MEM[32650] + MEM[32685];
assign MEM[40941] = MEM[32654] + MEM[32669];
assign MEM[40942] = MEM[32657] + MEM[32766];
assign MEM[40943] = MEM[32660] + MEM[32663];
assign MEM[40944] = MEM[32662] + MEM[32702];
assign MEM[40945] = MEM[32663] + MEM[32782];
assign MEM[40946] = MEM[32666] + MEM[32671];
assign MEM[40947] = MEM[32667] + MEM[32713];
assign MEM[40948] = MEM[32668] + MEM[32711];
assign MEM[40949] = MEM[32669] + MEM[32738];
assign MEM[40950] = MEM[32671] + MEM[32729];
assign MEM[40951] = MEM[32673] + MEM[32768];
assign MEM[40952] = MEM[32673] + MEM[32851];
assign MEM[40953] = MEM[32674] + MEM[32700];
assign MEM[40954] = MEM[32675] + MEM[32737];
assign MEM[40955] = MEM[32675] + MEM[32782];
assign MEM[40956] = MEM[32677] + MEM[32694];
assign MEM[40957] = MEM[32680] + MEM[32727];
assign MEM[40958] = MEM[32680] + MEM[32887];
assign MEM[40959] = MEM[32681] + MEM[32707];
assign MEM[40960] = MEM[32682] + MEM[32805];
assign MEM[40961] = MEM[32687] + MEM[32694];
assign MEM[40962] = MEM[32687] + MEM[32723];
assign MEM[40963] = MEM[32688] + MEM[32735];
assign MEM[40964] = MEM[32688] + MEM[32776];
assign MEM[40965] = MEM[32697] + MEM[32734];
assign MEM[40966] = MEM[32697] + MEM[32810];
assign MEM[40967] = MEM[32710] + MEM[32819];
assign MEM[40968] = MEM[32710] + MEM[32870];
assign MEM[40969] = MEM[32711] + MEM[32936];
assign MEM[40970] = MEM[32712] + MEM[32731];
assign MEM[40971] = MEM[32712] + MEM[32743];
assign MEM[40972] = MEM[32713] + MEM[32756];
assign MEM[40973] = MEM[32717] + MEM[32836];
assign MEM[40974] = MEM[32718] + MEM[32727];
assign MEM[40975] = MEM[32718] + MEM[32730];
assign MEM[40976] = MEM[32719] + MEM[32915];
assign MEM[40977] = MEM[32723] + MEM[32824];
assign MEM[40978] = MEM[32730] + MEM[32831];
assign MEM[40979] = MEM[32731] + MEM[32869];
assign MEM[40980] = MEM[32733] + MEM[32853];
assign MEM[40981] = MEM[32734] + MEM[32768];
assign MEM[40982] = MEM[32735] + MEM[32752];
assign MEM[40983] = MEM[32737] + MEM[32798];
assign MEM[40984] = MEM[32739] + MEM[32741];
assign MEM[40985] = MEM[32739] + MEM[32878];
assign MEM[40986] = MEM[32741] + MEM[32872];
assign MEM[40987] = MEM[32743] + MEM[32750];
assign MEM[40988] = MEM[32750] + MEM[32861];
assign MEM[40989] = MEM[32752] + MEM[32756];
assign MEM[40990] = MEM[32754] + MEM[32763];
assign MEM[40991] = MEM[32754] + MEM[32940];
assign MEM[40992] = MEM[32755] + MEM[32778];
assign MEM[40993] = MEM[32755] + MEM[32839];
assign MEM[40994] = MEM[32757] + MEM[32819];
assign MEM[40995] = MEM[32757] + MEM[32899];
assign MEM[40996] = MEM[32759] + MEM[32813];
assign MEM[40997] = MEM[32759] + MEM[32885];
assign MEM[40998] = MEM[32760] + MEM[32776];
assign MEM[40999] = MEM[32760] + MEM[32889];
assign MEM[41000] = MEM[32764] + MEM[32931];
assign MEM[41001] = MEM[32764] + MEM[32939];
assign MEM[41002] = MEM[32766] + MEM[32959];
assign MEM[41003] = MEM[32777] + MEM[32830];
assign MEM[41004] = MEM[32777] + MEM[32964];
assign MEM[41005] = MEM[32778] + MEM[32883];
assign MEM[41006] = MEM[32786] + MEM[32799];
assign MEM[41007] = MEM[32786] + MEM[32845];
assign MEM[41008] = MEM[32787] + MEM[32808];
assign MEM[41009] = MEM[32787] + MEM[32844];
assign MEM[41010] = MEM[32789] + MEM[32805];
assign MEM[41011] = MEM[32789] + MEM[32823];
assign MEM[41012] = MEM[32790] + MEM[33030];
assign MEM[41013] = MEM[32790] + MEM[33157];
assign MEM[41014] = MEM[32799] + MEM[32881];
assign MEM[41015] = MEM[32808] + MEM[32964];
assign MEM[41016] = MEM[32810] + MEM[32824];
assign MEM[41017] = MEM[32813] + MEM[32821];
assign MEM[41018] = MEM[32821] + MEM[32912];
assign MEM[41019] = MEM[32823] + MEM[32869];
assign MEM[41020] = MEM[32830] + MEM[32871];
assign MEM[41021] = MEM[32831] + MEM[32860];
assign MEM[41022] = MEM[32835] + MEM[32856];
assign MEM[41023] = MEM[32835] + MEM[32868];
assign MEM[41024] = MEM[32836] + MEM[32879];
assign MEM[41025] = MEM[32839] + MEM[32844];
assign MEM[41026] = MEM[32845] + MEM[32856];
assign MEM[41027] = MEM[32846] + MEM[32857];
assign MEM[41028] = MEM[32846] + MEM[32907];
assign MEM[41029] = MEM[32847] + MEM[32871];
assign MEM[41030] = MEM[32847] + MEM[32878];
assign MEM[41031] = MEM[32849] + MEM[32946];
assign MEM[41032] = MEM[32849] + MEM[33016];
assign MEM[41033] = MEM[32851] + MEM[32879];
assign MEM[41034] = MEM[32852] + MEM[32861];
assign MEM[41035] = MEM[32852] + MEM[33050];
assign MEM[41036] = MEM[32853] + MEM[32952];
assign MEM[41037] = MEM[32854] + MEM[32889];
assign MEM[41038] = MEM[32854] + MEM[32916];
assign MEM[41039] = MEM[32857] + MEM[32874];
assign MEM[41040] = MEM[32860] + MEM[32919];
assign MEM[41041] = MEM[32866] + MEM[32916];
assign MEM[41042] = MEM[32866] + MEM[32934];
assign MEM[41043] = MEM[32868] + MEM[32937];
assign MEM[41044] = MEM[32870] + MEM[32980];
assign MEM[41045] = MEM[32872] + MEM[32951];
assign MEM[41046] = MEM[32874] + MEM[32907];
assign MEM[41047] = MEM[32881] + MEM[32952];
assign MEM[41048] = MEM[32883] + MEM[32899];
assign MEM[41049] = MEM[32885] + MEM[33011];
assign MEM[41050] = MEM[32886] + MEM[32887];
assign MEM[41051] = MEM[32886] + MEM[32895];
assign MEM[41052] = MEM[32895] + MEM[32960];
assign MEM[41053] = MEM[32903] + MEM[32927];
assign MEM[41054] = MEM[32903] + MEM[33024];
assign MEM[41055] = MEM[32905] + MEM[32915];
assign MEM[41056] = MEM[32905] + MEM[32962];
assign MEM[41057] = MEM[32911] + MEM[32955];
assign MEM[41058] = MEM[32911] + MEM[32962];
assign MEM[41059] = MEM[32912] + MEM[33084];
assign MEM[41060] = MEM[32919] + MEM[32996];
assign MEM[41061] = MEM[32922] + MEM[32926];
assign MEM[41062] = MEM[32922] + MEM[32993];
assign MEM[41063] = MEM[32923] + MEM[32939];
assign MEM[41064] = MEM[32923] + MEM[33105];
assign MEM[41065] = MEM[32926] + MEM[33093];
assign MEM[41066] = MEM[32927] + MEM[33030];
assign MEM[41067] = MEM[32931] + MEM[32967];
assign MEM[41068] = MEM[32932] + MEM[32960];
assign MEM[41069] = MEM[32932] + MEM[33022];
assign MEM[41070] = MEM[32933] + MEM[32934];
assign MEM[41071] = MEM[32933] + MEM[32947];
assign MEM[41072] = MEM[32936] + MEM[33066];
assign MEM[41073] = MEM[32937] + MEM[32993];
assign MEM[41074] = MEM[32940] + MEM[32996];
assign MEM[41075] = MEM[32943] + MEM[32947];
assign MEM[41076] = MEM[32943] + MEM[33081];
assign MEM[41077] = MEM[32945] + MEM[32965];
assign MEM[41078] = MEM[32945] + MEM[32998];
assign MEM[41079] = MEM[32946] + MEM[32983];
assign MEM[41080] = MEM[32950] + MEM[33010];
assign MEM[41081] = MEM[32950] + MEM[33066];
assign MEM[41082] = MEM[32951] + MEM[33007];
assign MEM[41083] = MEM[32954] + MEM[33018];
assign MEM[41084] = MEM[32955] + MEM[33048];
assign MEM[41085] = MEM[32957] + MEM[32987];
assign MEM[41086] = MEM[32957] + MEM[33017];
assign MEM[41087] = MEM[32959] + MEM[32998];
assign MEM[41088] = MEM[32965] + MEM[33057];
assign MEM[41089] = MEM[32966] + MEM[33072];
assign MEM[41090] = MEM[32966] + MEM[33103];
assign MEM[41091] = MEM[32967] + MEM[32986];
assign MEM[41092] = MEM[32972] + MEM[32973];
assign MEM[41093] = MEM[32972] + MEM[33008];
assign MEM[41094] = MEM[32973] + MEM[33109];
assign MEM[41095] = MEM[32975] + MEM[33019];
assign MEM[41096] = MEM[32975] + MEM[33077];
assign MEM[41097] = MEM[32978] + MEM[32980];
assign MEM[41098] = MEM[32978] + MEM[33064];
assign MEM[41099] = MEM[32983] + MEM[32987];
assign MEM[41100] = MEM[32984] + MEM[33009];
assign MEM[41101] = MEM[32984] + MEM[33207];
assign MEM[41102] = MEM[32986] + MEM[33017];
assign MEM[41103] = MEM[32997] + MEM[33010];
assign MEM[41104] = MEM[32997] + MEM[33162];
assign MEM[41105] = MEM[32999] + MEM[33019];
assign MEM[41106] = MEM[32999] + MEM[33028];
assign MEM[41107] = MEM[33006] + MEM[33049];
assign MEM[41108] = MEM[33006] + MEM[33054];
assign MEM[41109] = MEM[33007] + MEM[33126];
assign MEM[41110] = MEM[33008] + MEM[33068];
assign MEM[41111] = MEM[33009] + MEM[33020];
assign MEM[41112] = MEM[33011] + MEM[33024];
assign MEM[41113] = MEM[33012] + MEM[33014];
assign MEM[41114] = MEM[33012] + MEM[33107];
assign MEM[41115] = MEM[33014] + MEM[33016];
assign MEM[41116] = MEM[33018] + MEM[33122];
assign MEM[41117] = MEM[33020] + MEM[33022];
assign MEM[41118] = MEM[33023] + MEM[33028];
assign MEM[41119] = MEM[33023] + MEM[33057];
assign MEM[41120] = MEM[33026] + MEM[33080];
assign MEM[41121] = MEM[33026] + MEM[33101];
assign MEM[41122] = MEM[33027] + MEM[33144];
assign MEM[41123] = MEM[33027] + MEM[33253];
assign MEM[41124] = MEM[33037] + MEM[33044];
assign MEM[41125] = MEM[33037] + MEM[33061];
assign MEM[41126] = MEM[33042] + MEM[33044];
assign MEM[41127] = MEM[33042] + MEM[33096];
assign MEM[41128] = MEM[33043] + MEM[33082];
assign MEM[41129] = MEM[33043] + MEM[33088];
assign MEM[41130] = MEM[33048] + MEM[33067];
assign MEM[41131] = MEM[33049] + MEM[33055];
assign MEM[41132] = MEM[33050] + MEM[33148];
assign MEM[41133] = MEM[33054] + MEM[33081];
assign MEM[41134] = MEM[33055] + MEM[33101];
assign MEM[41135] = MEM[33061] + MEM[33156];
assign MEM[41136] = MEM[33062] + MEM[33079];
assign MEM[41137] = MEM[33062] + MEM[33088];
assign MEM[41138] = MEM[33063] + MEM[33120];
assign MEM[41139] = MEM[33063] + MEM[33140];
assign MEM[41140] = MEM[33064] + MEM[33111];
assign MEM[41141] = MEM[33067] + MEM[33124];
assign MEM[41142] = MEM[33068] + MEM[33069];
assign MEM[41143] = MEM[33069] + MEM[33078];
assign MEM[41144] = MEM[33070] + MEM[33117];
assign MEM[41145] = MEM[33070] + MEM[33135];
assign MEM[41146] = MEM[33072] + MEM[33114];
assign MEM[41147] = MEM[33073] + MEM[33080];
assign MEM[41148] = MEM[33073] + MEM[33104];
assign MEM[41149] = MEM[33077] + MEM[33214];
assign MEM[41150] = MEM[33078] + MEM[33220];
assign MEM[41151] = MEM[33079] + MEM[33141];
assign MEM[41152] = MEM[33082] + MEM[33224];
assign MEM[41153] = MEM[33084] + MEM[33131];
assign MEM[41154] = MEM[33086] + MEM[33092];
assign MEM[41155] = MEM[33086] + MEM[33093];
assign MEM[41156] = MEM[33087] + MEM[33104];
assign MEM[41157] = MEM[33087] + MEM[33109];
assign MEM[41158] = MEM[33092] + MEM[33110];
assign MEM[41159] = MEM[33096] + MEM[33159];
assign MEM[41160] = MEM[33097] + MEM[33133];
assign MEM[41161] = MEM[33097] + MEM[33150];
assign MEM[41162] = MEM[33103] + MEM[33108];
assign MEM[41163] = MEM[33105] + MEM[33153];
assign MEM[41164] = MEM[33107] + MEM[33138];
assign MEM[41165] = MEM[33108] + MEM[33166];
assign MEM[41166] = MEM[33110] + MEM[33112];
assign MEM[41167] = MEM[33111] + MEM[33127];
assign MEM[41168] = MEM[33112] + MEM[33115];
assign MEM[41169] = MEM[33114] + MEM[33215];
assign MEM[41170] = MEM[33115] + MEM[33119];
assign MEM[41171] = MEM[33116] + MEM[33131];
assign MEM[41172] = MEM[33116] + MEM[33162];
assign MEM[41173] = MEM[33117] + MEM[33153];
assign MEM[41174] = MEM[33118] + MEM[33119];
assign MEM[41175] = MEM[33118] + MEM[33149];
assign MEM[41176] = MEM[33120] + MEM[33130];
assign MEM[41177] = MEM[33122] + MEM[33176];
assign MEM[41178] = MEM[33124] + MEM[33156];
assign MEM[41179] = MEM[33125] + MEM[33137];
assign MEM[41180] = MEM[33125] + MEM[33154];
assign MEM[41181] = MEM[33126] + MEM[33178];
assign MEM[41182] = MEM[33127] + MEM[33144];
assign MEM[41183] = MEM[33128] + MEM[33159];
assign MEM[41184] = MEM[33128] + MEM[33178];
assign MEM[41185] = MEM[33129] + MEM[33145];
assign MEM[41186] = MEM[33129] + MEM[33146];
assign MEM[41187] = MEM[33130] + MEM[33170];
assign MEM[41188] = MEM[33132] + MEM[33167];
assign MEM[41189] = MEM[33132] + MEM[33184];
assign MEM[41190] = MEM[33133] + MEM[33158];
assign MEM[41191] = MEM[33135] + MEM[33158];
assign MEM[41192] = MEM[33137] + MEM[33262];
assign MEM[41193] = MEM[33138] + MEM[33224];
assign MEM[41194] = MEM[33139] + MEM[33141];
assign MEM[41195] = MEM[33139] + MEM[33229];
assign MEM[41196] = MEM[33140] + MEM[33176];
assign MEM[41197] = MEM[33143] + MEM[33177];
assign MEM[41198] = MEM[33143] + MEM[33201];
assign MEM[41199] = MEM[33145] + MEM[33161];
assign MEM[41200] = MEM[33146] + MEM[33225];
assign MEM[41201] = MEM[33147] + MEM[33148];
assign MEM[41202] = MEM[33147] + MEM[33161];
assign MEM[41203] = MEM[33149] + MEM[33298];
assign MEM[41204] = MEM[33150] + MEM[33164];
assign MEM[41205] = MEM[33152] + MEM[33157];
assign MEM[41206] = MEM[33152] + MEM[33192];
assign MEM[41207] = MEM[33154] + MEM[33196];
assign MEM[41208] = MEM[33160] + MEM[33172];
assign MEM[41209] = MEM[33160] + MEM[33203];
assign MEM[41210] = MEM[33164] + MEM[33226];
assign MEM[41211] = MEM[33165] + MEM[33183];
assign MEM[41212] = MEM[33165] + MEM[33218];
assign MEM[41213] = MEM[33166] + MEM[33214];
assign MEM[41214] = MEM[33167] + MEM[33173];
assign MEM[41215] = MEM[33170] + MEM[33171];
assign MEM[41216] = MEM[33171] + MEM[33241];
assign MEM[41217] = MEM[33172] + MEM[33261];
assign MEM[41218] = MEM[33173] + MEM[33181];
assign MEM[41219] = MEM[33174] + MEM[33247];
assign MEM[41220] = MEM[33174] + MEM[33273];
assign MEM[41221] = MEM[33175] + MEM[33188];
assign MEM[41222] = MEM[33175] + MEM[33267];
assign MEM[41223] = MEM[33177] + MEM[33206];
assign MEM[41224] = MEM[33179] + MEM[33192];
assign MEM[41225] = MEM[33179] + MEM[33208];
assign MEM[41226] = MEM[33181] + MEM[33183];
assign MEM[41227] = MEM[33182] + MEM[33198];
assign MEM[41228] = MEM[33182] + MEM[33215];
assign MEM[41229] = MEM[33184] + MEM[33202];
assign MEM[41230] = MEM[33186] + MEM[33193];
assign MEM[41231] = MEM[33186] + MEM[33245];
assign MEM[41232] = MEM[33187] + MEM[33189];
assign MEM[41233] = MEM[33187] + MEM[33292];
assign MEM[41234] = MEM[33188] + MEM[33190];
assign MEM[41235] = MEM[33189] + MEM[33237];
assign MEM[41236] = MEM[33190] + MEM[33246];
assign MEM[41237] = MEM[33193] + MEM[33196];
assign MEM[41238] = MEM[33198] + MEM[33255];
assign MEM[41239] = MEM[33200] + MEM[33211];
assign MEM[41240] = MEM[33200] + MEM[33221];
assign MEM[41241] = MEM[33201] + MEM[33238];
assign MEM[41242] = MEM[33202] + MEM[33263];
assign MEM[41243] = MEM[33203] + MEM[33248];
assign MEM[41244] = MEM[33205] + MEM[33217];
assign MEM[41245] = MEM[33205] + MEM[33231];
assign MEM[41246] = MEM[33206] + MEM[33219];
assign MEM[41247] = MEM[33207] + MEM[33313];
assign MEM[41248] = MEM[33208] + MEM[33256];
assign MEM[41249] = MEM[33211] + MEM[33242];
assign MEM[41250] = MEM[33212] + MEM[33213];
assign MEM[41251] = MEM[33212] + MEM[33265];
assign MEM[41252] = MEM[33213] + MEM[33294];
assign MEM[41253] = MEM[33216] + MEM[33231];
assign MEM[41254] = MEM[33216] + MEM[33234];
assign MEM[41255] = MEM[33217] + MEM[33295];
assign MEM[41256] = MEM[33218] + MEM[33225];
assign MEM[41257] = MEM[33219] + MEM[33248];
assign MEM[41258] = MEM[33220] + MEM[33288];
assign MEM[41259] = MEM[33221] + MEM[33250];
assign MEM[41260] = MEM[33223] + MEM[33233];
assign MEM[41261] = MEM[33223] + MEM[33244];
assign MEM[41262] = MEM[33226] + MEM[33240];
assign MEM[41263] = MEM[33229] + MEM[33353];
assign MEM[41264] = MEM[33230] + MEM[33305];
assign MEM[41265] = MEM[33230] + MEM[33307];
assign MEM[41266] = MEM[33232] + MEM[33245];
assign MEM[41267] = MEM[33232] + MEM[33261];
assign MEM[41268] = MEM[33233] + MEM[33258];
assign MEM[41269] = MEM[33234] + MEM[33387];
assign MEM[41270] = MEM[33236] + MEM[33259];
assign MEM[41271] = MEM[33236] + MEM[33264];
assign MEM[41272] = MEM[33237] + MEM[33265];
assign MEM[41273] = MEM[33238] + MEM[33240];
assign MEM[41274] = MEM[33241] + MEM[33269];
assign MEM[41275] = MEM[33242] + MEM[33340];
assign MEM[41276] = MEM[33244] + MEM[33275];
assign MEM[41277] = MEM[33246] + MEM[33253];
assign MEM[41278] = MEM[33247] + MEM[33308];
assign MEM[41279] = MEM[33249] + MEM[33289];
assign MEM[41280] = MEM[33249] + MEM[33302];
assign MEM[41281] = MEM[33250] + MEM[33317];
assign MEM[41282] = MEM[33251] + MEM[33267];
assign MEM[41283] = MEM[33251] + MEM[33285];
assign MEM[41284] = MEM[33254] + MEM[33288];
assign MEM[41285] = MEM[33254] + MEM[33298];
assign MEM[41286] = MEM[33255] + MEM[33299];
assign MEM[41287] = MEM[33256] + MEM[33260];
assign MEM[41288] = MEM[33258] + MEM[33291];
assign MEM[41289] = MEM[33259] + MEM[33323];
assign MEM[41290] = MEM[33260] + MEM[33280];
assign MEM[41291] = MEM[33262] + MEM[33299];
assign MEM[41292] = MEM[33263] + MEM[33279];
assign MEM[41293] = MEM[33264] + MEM[33266];
assign MEM[41294] = MEM[33266] + MEM[33323];
assign MEM[41295] = MEM[33268] + MEM[33269];
assign MEM[41296] = MEM[33268] + MEM[33338];
assign MEM[41297] = MEM[33270] + MEM[33271];
assign MEM[41298] = MEM[33270] + MEM[33278];
assign MEM[41299] = MEM[33271] + MEM[33292];
assign MEM[41300] = MEM[33272] + MEM[33274];
assign MEM[41301] = MEM[33272] + MEM[33321];
assign MEM[41302] = MEM[33273] + MEM[33321];
assign MEM[41303] = MEM[33274] + MEM[33275];
assign MEM[41304] = MEM[33276] + MEM[33281];
assign MEM[41305] = MEM[33276] + MEM[33312];
assign MEM[41306] = MEM[33277] + MEM[33294];
assign MEM[41307] = MEM[33277] + MEM[33333];
assign MEM[41308] = MEM[33278] + MEM[33325];
assign MEM[41309] = MEM[33279] + MEM[33302];
assign MEM[41310] = MEM[33280] + MEM[33284];
assign MEM[41311] = MEM[33281] + MEM[33368];
assign MEM[41312] = MEM[33284] + MEM[33295];
assign MEM[41313] = MEM[33285] + MEM[33310];
assign MEM[41314] = MEM[33286] + MEM[33311];
assign MEM[41315] = MEM[33286] + MEM[33433];
assign MEM[41316] = MEM[33287] + MEM[33320];
assign MEM[41317] = MEM[33287] + MEM[33375];
assign MEM[41318] = MEM[33289] + MEM[33316];
assign MEM[41319] = MEM[33290] + MEM[33291];
assign MEM[41320] = MEM[33290] + MEM[33297];
assign MEM[41321] = MEM[33293] + MEM[33297];
assign MEM[41322] = MEM[33293] + MEM[33320];
assign MEM[41323] = MEM[33296] + MEM[33322];
assign MEM[41324] = MEM[33296] + MEM[33337];
assign MEM[41325] = MEM[33300] + MEM[33310];
assign MEM[41326] = MEM[33300] + MEM[33325];
assign MEM[41327] = MEM[33304] + MEM[33314];
assign MEM[41328] = MEM[33304] + MEM[33336];
assign MEM[41329] = MEM[33305] + MEM[33309];
assign MEM[41330] = MEM[33307] + MEM[33324];
assign MEM[41331] = MEM[33308] + MEM[33552];
assign MEM[41332] = MEM[33309] + MEM[33341];
assign MEM[41333] = MEM[33311] + MEM[33333];
assign MEM[41334] = MEM[33312] + MEM[33364];
assign MEM[41335] = MEM[33313] + MEM[33367];
assign MEM[41336] = MEM[33314] + MEM[33358];
assign MEM[41337] = MEM[33315] + MEM[33334];
assign MEM[41338] = MEM[33315] + MEM[33380];
assign MEM[41339] = MEM[33316] + MEM[33384];
assign MEM[41340] = MEM[33317] + MEM[33327];
assign MEM[41341] = MEM[33318] + MEM[33363];
assign MEM[41342] = MEM[33318] + MEM[33443];
assign MEM[41343] = MEM[33322] + MEM[33332];
assign MEM[41344] = MEM[33324] + MEM[33341];
assign MEM[41345] = MEM[33326] + MEM[33346];
assign MEM[41346] = MEM[33326] + MEM[33348];
assign MEM[41347] = MEM[33327] + MEM[33332];
assign MEM[41348] = MEM[33329] + MEM[33330];
assign MEM[41349] = MEM[33329] + MEM[33431];
assign MEM[41350] = MEM[33330] + MEM[33455];
assign MEM[41351] = MEM[33331] + MEM[33360];
assign MEM[41352] = MEM[33331] + MEM[33402];
assign MEM[41353] = MEM[33334] + MEM[33379];
assign MEM[41354] = MEM[33335] + MEM[33354];
assign MEM[41355] = MEM[33335] + MEM[33373];
assign MEM[41356] = MEM[33336] + MEM[33371];
assign MEM[41357] = MEM[33337] + MEM[33352];
assign MEM[41358] = MEM[33338] + MEM[33419];
assign MEM[41359] = MEM[33339] + MEM[33343];
assign MEM[41360] = MEM[33339] + MEM[33362];
assign MEM[41361] = MEM[33340] + MEM[33352];
assign MEM[41362] = MEM[33343] + MEM[33344];
assign MEM[41363] = MEM[33344] + MEM[33543];
assign MEM[41364] = MEM[33346] + MEM[33388];
assign MEM[41365] = MEM[33347] + MEM[33356];
assign MEM[41366] = MEM[33347] + MEM[33400];
assign MEM[41367] = MEM[33348] + MEM[33357];
assign MEM[41368] = MEM[33350] + MEM[33412];
assign MEM[41369] = MEM[33350] + MEM[33491];
assign MEM[41370] = MEM[33351] + MEM[33355];
assign MEM[41371] = MEM[33351] + MEM[33374];
assign MEM[41372] = MEM[33353] + MEM[33439];
assign MEM[41373] = MEM[33354] + MEM[33360];
assign MEM[41374] = MEM[33355] + MEM[33359];
assign MEM[41375] = MEM[33356] + MEM[33361];
assign MEM[41376] = MEM[33357] + MEM[33359];
assign MEM[41377] = MEM[33358] + MEM[33429];
assign MEM[41378] = MEM[33361] + MEM[33378];
assign MEM[41379] = MEM[33362] + MEM[33413];
assign MEM[41380] = MEM[33363] + MEM[33400];
assign MEM[41381] = MEM[33364] + MEM[33378];
assign MEM[41382] = MEM[33366] + MEM[33367];
assign MEM[41383] = MEM[33366] + MEM[33373];
assign MEM[41384] = MEM[33368] + MEM[33406];
assign MEM[41385] = MEM[33370] + MEM[33379];
assign MEM[41386] = MEM[33370] + MEM[33390];
assign MEM[41387] = MEM[33371] + MEM[33478];
assign MEM[41388] = MEM[33374] + MEM[33377];
assign MEM[41389] = MEM[33375] + MEM[33401];
assign MEM[41390] = MEM[33377] + MEM[33444];
assign MEM[41391] = MEM[33380] + MEM[33385];
assign MEM[41392] = MEM[33381] + MEM[33392];
assign MEM[41393] = MEM[33381] + MEM[33413];
assign MEM[41394] = MEM[33382] + MEM[33432];
assign MEM[41395] = MEM[33382] + MEM[33450];
assign MEM[41396] = MEM[33383] + MEM[33410];
assign MEM[41397] = MEM[33383] + MEM[33431];
assign MEM[41398] = MEM[33384] + MEM[33403];
assign MEM[41399] = MEM[33385] + MEM[33434];
assign MEM[41400] = MEM[33386] + MEM[33388];
assign MEM[41401] = MEM[33386] + MEM[33411];
assign MEM[41402] = MEM[33387] + MEM[33463];
assign MEM[41403] = MEM[33390] + MEM[33408];
assign MEM[41404] = MEM[33391] + MEM[33395];
assign MEM[41405] = MEM[33391] + MEM[33420];
assign MEM[41406] = MEM[33392] + MEM[33475];
assign MEM[41407] = MEM[33393] + MEM[33403];
assign MEM[41408] = MEM[33393] + MEM[33417];
assign MEM[41409] = MEM[33394] + MEM[33398];
assign MEM[41410] = MEM[33394] + MEM[33406];
assign MEM[41411] = MEM[33395] + MEM[33440];
assign MEM[41412] = MEM[33396] + MEM[33419];
assign MEM[41413] = MEM[33396] + MEM[33446];
assign MEM[41414] = MEM[33398] + MEM[33424];
assign MEM[41415] = MEM[33399] + MEM[33412];
assign MEM[41416] = MEM[33399] + MEM[33418];
assign MEM[41417] = MEM[33401] + MEM[33482];
assign MEM[41418] = MEM[33402] + MEM[33410];
assign MEM[41419] = MEM[33405] + MEM[33423];
assign MEM[41420] = MEM[33405] + MEM[33437];
assign MEM[41421] = MEM[33407] + MEM[33409];
assign MEM[41422] = MEM[33407] + MEM[33418];
assign MEM[41423] = MEM[33408] + MEM[33488];
assign MEM[41424] = MEM[33409] + MEM[33571];
assign MEM[41425] = MEM[33411] + MEM[33451];
assign MEM[41426] = MEM[33416] + MEM[33420];
assign MEM[41427] = MEM[33416] + MEM[33586];
assign MEM[41428] = MEM[33417] + MEM[33422];
assign MEM[41429] = MEM[33422] + MEM[33442];
assign MEM[41430] = MEM[33423] + MEM[33435];
assign MEM[41431] = MEM[33424] + MEM[33428];
assign MEM[41432] = MEM[33425] + MEM[33437];
assign MEM[41433] = MEM[33425] + MEM[33438];
assign MEM[41434] = MEM[33428] + MEM[33443];
assign MEM[41435] = MEM[33429] + MEM[33494];
assign MEM[41436] = MEM[33430] + MEM[33458];
assign MEM[41437] = MEM[33430] + MEM[33465];
assign MEM[41438] = MEM[33432] + MEM[33501];
assign MEM[41439] = MEM[33433] + MEM[33468];
assign MEM[41440] = MEM[33434] + MEM[33464];
assign MEM[41441] = MEM[33435] + MEM[33529];
assign MEM[41442] = MEM[33436] + MEM[33455];
assign MEM[41443] = MEM[33436] + MEM[33471];
assign MEM[41444] = MEM[33438] + MEM[33446];
assign MEM[41445] = MEM[33439] + MEM[33449];
assign MEM[41446] = MEM[33440] + MEM[33537];
assign MEM[41447] = MEM[33441] + MEM[33451];
assign MEM[41448] = MEM[33441] + MEM[33460];
assign MEM[41449] = MEM[33442] + MEM[33452];
assign MEM[41450] = MEM[33444] + MEM[33453];
assign MEM[41451] = MEM[33445] + MEM[33449];
assign MEM[41452] = MEM[33445] + MEM[33547];
assign MEM[41453] = MEM[33448] + MEM[33457];
assign MEM[41454] = MEM[33448] + MEM[33532];
assign MEM[41455] = MEM[33450] + MEM[33478];
assign MEM[41456] = MEM[33452] + MEM[33548];
assign MEM[41457] = MEM[33453] + MEM[33482];
assign MEM[41458] = MEM[33456] + MEM[33495];
assign MEM[41459] = MEM[33456] + MEM[33583];
assign MEM[41460] = MEM[33457] + MEM[33458];
assign MEM[41461] = MEM[33459] + MEM[33491];
assign MEM[41462] = MEM[33459] + MEM[33511];
assign MEM[41463] = MEM[33460] + MEM[33502];
assign MEM[41464] = MEM[33461] + MEM[33485];
assign MEM[41465] = MEM[33461] + MEM[33496];
assign MEM[41466] = MEM[33463] + MEM[33473];
assign MEM[41467] = MEM[33464] + MEM[33556];
assign MEM[41468] = MEM[33465] + MEM[33496];
assign MEM[41469] = MEM[33466] + MEM[33468];
assign MEM[41470] = MEM[33466] + MEM[33503];
assign MEM[41471] = MEM[33467] + MEM[33492];
assign MEM[41472] = MEM[33467] + MEM[33507];
assign MEM[41473] = MEM[33469] + MEM[33488];
assign MEM[41474] = MEM[33469] + MEM[33570];
assign MEM[41475] = MEM[33471] + MEM[33486];
assign MEM[41476] = MEM[33472] + MEM[33477];
assign MEM[41477] = MEM[33472] + MEM[33537];
assign MEM[41478] = MEM[33473] + MEM[33516];
assign MEM[41479] = MEM[33475] + MEM[33504];
assign MEM[41480] = MEM[33477] + MEM[33487];
assign MEM[41481] = MEM[33479] + MEM[33480];
assign MEM[41482] = MEM[33479] + MEM[33526];
assign MEM[41483] = MEM[33480] + MEM[33504];
assign MEM[41484] = MEM[33481] + MEM[33493];
assign MEM[41485] = MEM[33481] + MEM[33513];
assign MEM[41486] = MEM[33484] + MEM[33508];
assign MEM[41487] = MEM[33484] + MEM[33565];
assign MEM[41488] = MEM[33485] + MEM[33487];
assign MEM[41489] = MEM[33486] + MEM[33506];
assign MEM[41490] = MEM[33489] + MEM[33494];
assign MEM[41491] = MEM[33489] + MEM[33571];
assign MEM[41492] = MEM[33492] + MEM[33535];
assign MEM[41493] = MEM[33493] + MEM[33523];
assign MEM[41494] = MEM[33495] + MEM[33506];
assign MEM[41495] = MEM[33497] + MEM[33500];
assign MEM[41496] = MEM[33497] + MEM[33501];
assign MEM[41497] = MEM[33498] + MEM[33515];
assign MEM[41498] = MEM[33498] + MEM[33541];
assign MEM[41499] = MEM[33500] + MEM[33514];
assign MEM[41500] = MEM[33502] + MEM[33587];
assign MEM[41501] = MEM[33503] + MEM[33513];
assign MEM[41502] = MEM[33505] + MEM[33535];
assign MEM[41503] = MEM[33505] + MEM[33565];
assign MEM[41504] = MEM[33507] + MEM[33536];
assign MEM[41505] = MEM[33508] + MEM[33689];
assign MEM[41506] = MEM[33509] + MEM[33517];
assign MEM[41507] = MEM[33509] + MEM[33521];
assign MEM[41508] = MEM[33510] + MEM[33540];
assign MEM[41509] = MEM[33510] + MEM[33597];
assign MEM[41510] = MEM[33511] + MEM[33514];
assign MEM[41511] = MEM[33515] + MEM[33519];
assign MEM[41512] = MEM[33516] + MEM[33578];
assign MEM[41513] = MEM[33517] + MEM[33560];
assign MEM[41514] = MEM[33518] + MEM[33527];
assign MEM[41515] = MEM[33518] + MEM[33584];
assign MEM[41516] = MEM[33519] + MEM[33525];
assign MEM[41517] = MEM[33520] + MEM[33526];
assign MEM[41518] = MEM[33520] + MEM[33528];
assign MEM[41519] = MEM[33521] + MEM[33539];
assign MEM[41520] = MEM[33522] + MEM[33534];
assign MEM[41521] = MEM[33522] + MEM[33635];
assign MEM[41522] = MEM[33523] + MEM[33562];
assign MEM[41523] = MEM[33525] + MEM[33527];
assign MEM[41524] = MEM[33528] + MEM[33530];
assign MEM[41525] = MEM[33529] + MEM[33543];
assign MEM[41526] = MEM[33530] + MEM[33601];
assign MEM[41527] = MEM[33532] + MEM[33707];
assign MEM[41528] = MEM[33534] + MEM[33557];
assign MEM[41529] = MEM[33536] + MEM[33551];
assign MEM[41530] = MEM[33538] + MEM[33567];
assign MEM[41531] = MEM[33538] + MEM[33621];
assign MEM[41532] = MEM[33539] + MEM[33606];
assign MEM[41533] = MEM[33540] + MEM[33558];
assign MEM[41534] = MEM[33541] + MEM[33545];
assign MEM[41535] = MEM[33544] + MEM[33577];
assign MEM[41536] = MEM[33544] + MEM[33583];
assign MEM[41537] = MEM[33545] + MEM[33684];
assign MEM[41538] = MEM[33546] + MEM[33606];
assign MEM[41539] = MEM[33546] + MEM[33608];
assign MEM[41540] = MEM[33547] + MEM[33622];
assign MEM[41541] = MEM[33548] + MEM[33587];
assign MEM[41542] = MEM[33549] + MEM[33568];
assign MEM[41543] = MEM[33549] + MEM[33579];
assign MEM[41544] = MEM[33551] + MEM[33575];
assign MEM[41545] = MEM[33552] + MEM[33555];
assign MEM[41546] = MEM[33554] + MEM[33567];
assign MEM[41547] = MEM[33554] + MEM[33585];
assign MEM[41548] = MEM[33555] + MEM[33642];
assign MEM[41549] = MEM[33556] + MEM[33581];
assign MEM[41550] = MEM[33557] + MEM[33595];
assign MEM[41551] = MEM[33558] + MEM[33564];
assign MEM[41552] = MEM[33559] + MEM[33561];
assign MEM[41553] = MEM[33559] + MEM[33566];
assign MEM[41554] = MEM[33560] + MEM[33593];
assign MEM[41555] = MEM[33561] + MEM[33590];
assign MEM[41556] = MEM[33562] + MEM[33647];
assign MEM[41557] = MEM[33564] + MEM[33600];
assign MEM[41558] = MEM[33566] + MEM[33572];
assign MEM[41559] = MEM[33568] + MEM[33594];
assign MEM[41560] = MEM[33569] + MEM[33577];
assign MEM[41561] = MEM[33569] + MEM[33615];
assign MEM[41562] = MEM[33570] + MEM[33590];
assign MEM[41563] = MEM[33572] + MEM[33588];
assign MEM[41564] = MEM[33575] + MEM[33588];
assign MEM[41565] = MEM[33576] + MEM[33581];
assign MEM[41566] = MEM[33576] + MEM[33585];
assign MEM[41567] = MEM[33578] + MEM[33602];
assign MEM[41568] = MEM[33579] + MEM[33607];
assign MEM[41569] = MEM[33580] + MEM[33625];
assign MEM[41570] = MEM[33580] + MEM[33668];
assign MEM[41571] = MEM[33582] + MEM[33605];
assign MEM[41572] = MEM[33582] + MEM[33632];
assign MEM[41573] = MEM[33584] + MEM[33633];
assign MEM[41574] = MEM[33586] + MEM[33616];
assign MEM[41575] = MEM[33589] + MEM[33604];
assign MEM[41576] = MEM[33589] + MEM[33622];
assign MEM[41577] = MEM[33592] + MEM[33614];
assign MEM[41578] = MEM[33592] + MEM[33674];
assign MEM[41579] = MEM[33593] + MEM[33611];
assign MEM[41580] = MEM[33594] + MEM[33603];
assign MEM[41581] = MEM[33595] + MEM[33673];
assign MEM[41582] = MEM[33596] + MEM[33607];
assign MEM[41583] = MEM[33596] + MEM[33654];
assign MEM[41584] = MEM[33597] + MEM[33605];
assign MEM[41585] = MEM[33600] + MEM[33617];
assign MEM[41586] = MEM[33601] + MEM[33618];
assign MEM[41587] = MEM[33602] + MEM[33604];
assign MEM[41588] = MEM[33603] + MEM[33641];
assign MEM[41589] = MEM[33608] + MEM[33630];
assign MEM[41590] = MEM[33609] + MEM[33623];
assign MEM[41591] = MEM[33609] + MEM[33646];
assign MEM[41592] = MEM[33610] + MEM[33620];
assign MEM[41593] = MEM[33610] + MEM[33630];
assign MEM[41594] = MEM[33611] + MEM[33639];
assign MEM[41595] = MEM[33613] + MEM[33644];
assign MEM[41596] = MEM[33613] + MEM[33651];
assign MEM[41597] = MEM[33614] + MEM[33628];
assign MEM[41598] = MEM[33615] + MEM[33655];
assign MEM[41599] = MEM[33616] + MEM[33639];
assign MEM[41600] = MEM[33617] + MEM[33646];
assign MEM[41601] = MEM[33618] + MEM[33621];
assign MEM[41602] = MEM[33619] + MEM[33623];
assign MEM[41603] = MEM[33619] + MEM[33640];
assign MEM[41604] = MEM[33620] + MEM[33676];
assign MEM[41605] = MEM[33624] + MEM[33625];
assign MEM[41606] = MEM[33624] + MEM[33710];
assign MEM[41607] = MEM[33627] + MEM[33631];
assign MEM[41608] = MEM[33627] + MEM[33667];
assign MEM[41609] = MEM[33628] + MEM[33669];
assign MEM[41610] = MEM[33629] + MEM[33631];
assign MEM[41611] = MEM[33629] + MEM[33679];
assign MEM[41612] = MEM[33632] + MEM[33687];
assign MEM[41613] = MEM[33633] + MEM[33643];
assign MEM[41614] = MEM[33634] + MEM[33635];
assign MEM[41615] = MEM[33634] + MEM[33656];
assign MEM[41616] = MEM[33636] + MEM[33640];
assign MEM[41617] = MEM[33636] + MEM[33717];
assign MEM[41618] = MEM[33637] + MEM[33653];
assign MEM[41619] = MEM[33637] + MEM[33658];
assign MEM[41620] = MEM[33638] + MEM[33659];
assign MEM[41621] = MEM[33638] + MEM[33704];
assign MEM[41622] = MEM[33641] + MEM[33652];
assign MEM[41623] = MEM[33642] + MEM[33677];
assign MEM[41624] = MEM[33643] + MEM[33650];
assign MEM[41625] = MEM[33644] + MEM[33685];
assign MEM[41626] = MEM[33647] + MEM[33745];
assign MEM[41627] = MEM[33648] + MEM[33677];
assign MEM[41628] = MEM[33648] + MEM[33693];
assign MEM[41629] = MEM[33649] + MEM[33682];
assign MEM[41630] = MEM[33649] + MEM[33693];
assign MEM[41631] = MEM[33650] + MEM[33760];
assign MEM[41632] = MEM[33651] + MEM[33699];
assign MEM[41633] = MEM[33652] + MEM[33654];
assign MEM[41634] = MEM[33653] + MEM[33685];
assign MEM[41635] = MEM[33655] + MEM[33694];
assign MEM[41636] = MEM[33656] + MEM[33664];
assign MEM[41637] = MEM[33658] + MEM[33719];
assign MEM[41638] = MEM[33659] + MEM[33664];
assign MEM[41639] = MEM[33661] + MEM[33665];
assign MEM[41640] = MEM[33661] + MEM[33666];
assign MEM[41641] = MEM[33662] + MEM[33678];
assign MEM[41642] = MEM[33662] + MEM[33683];
assign MEM[41643] = MEM[33663] + MEM[33680];
assign MEM[41644] = MEM[33663] + MEM[33682];
assign MEM[41645] = MEM[33665] + MEM[33789];
assign MEM[41646] = MEM[33666] + MEM[33675];
assign MEM[41647] = MEM[33667] + MEM[33777];
assign MEM[41648] = MEM[33668] + MEM[33750];
assign MEM[41649] = MEM[33669] + MEM[33679];
assign MEM[41650] = MEM[33670] + MEM[33674];
assign MEM[41651] = MEM[33670] + MEM[33675];
assign MEM[41652] = MEM[33671] + MEM[33698];
assign MEM[41653] = MEM[33671] + MEM[33724];
assign MEM[41654] = MEM[33672] + MEM[33676];
assign MEM[41655] = MEM[33672] + MEM[33749];
assign MEM[41656] = MEM[33673] + MEM[33694];
assign MEM[41657] = MEM[33678] + MEM[33684];
assign MEM[41658] = MEM[33680] + MEM[33702];
assign MEM[41659] = MEM[33683] + MEM[33770];
assign MEM[41660] = MEM[33687] + MEM[33699];
assign MEM[41661] = MEM[33688] + MEM[33702];
assign MEM[41662] = MEM[33688] + MEM[33770];
assign MEM[41663] = MEM[33689] + MEM[33724];
assign MEM[41664] = MEM[33690] + MEM[33695];
assign MEM[41665] = MEM[33690] + MEM[33762];
assign MEM[41666] = MEM[33691] + MEM[33738];
assign MEM[41667] = MEM[33691] + MEM[33766];
assign MEM[41668] = MEM[33692] + MEM[33726];
assign MEM[41669] = MEM[33692] + MEM[33765];
assign MEM[41670] = MEM[33695] + MEM[33841];
assign MEM[41671] = MEM[33697] + MEM[33700];
assign MEM[41672] = MEM[33697] + MEM[33715];
assign MEM[41673] = MEM[33698] + MEM[33705];
assign MEM[41674] = MEM[33700] + MEM[33703];
assign MEM[41675] = MEM[33701] + MEM[33722];
assign MEM[41676] = MEM[33701] + MEM[33762];
assign MEM[41677] = MEM[33703] + MEM[33706];
assign MEM[41678] = MEM[33704] + MEM[33733];
assign MEM[41679] = MEM[33705] + MEM[33727];
assign MEM[41680] = MEM[33706] + MEM[33709];
assign MEM[41681] = MEM[33707] + MEM[33717];
assign MEM[41682] = MEM[33708] + MEM[33748];
assign MEM[41683] = MEM[33708] + MEM[33763];
assign MEM[41684] = MEM[33709] + MEM[33798];
assign MEM[41685] = MEM[33710] + MEM[33746];
assign MEM[41686] = MEM[33711] + MEM[33720];
assign MEM[41687] = MEM[33711] + MEM[33731];
assign MEM[41688] = MEM[33712] + MEM[33719];
assign MEM[41689] = MEM[33712] + MEM[33732];
assign MEM[41690] = MEM[33713] + MEM[33718];
assign MEM[41691] = MEM[33713] + MEM[33727];
assign MEM[41692] = MEM[33714] + MEM[33716];
assign MEM[41693] = MEM[33714] + MEM[33765];
assign MEM[41694] = MEM[33715] + MEM[33812];
assign MEM[41695] = MEM[33716] + MEM[33728];
assign MEM[41696] = MEM[33718] + MEM[33731];
assign MEM[41697] = MEM[33720] + MEM[33729];
assign MEM[41698] = MEM[33721] + MEM[33734];
assign MEM[41699] = MEM[33721] + MEM[33763];
assign MEM[41700] = MEM[33722] + MEM[33759];
assign MEM[41701] = MEM[33723] + MEM[33761];
assign MEM[41702] = MEM[33723] + MEM[33775];
assign MEM[41703] = MEM[33725] + MEM[33732];
assign MEM[41704] = MEM[33725] + MEM[33735];
assign MEM[41705] = MEM[33726] + MEM[33741];
assign MEM[41706] = MEM[33728] + MEM[33787];
assign MEM[41707] = MEM[33729] + MEM[33750];
assign MEM[41708] = MEM[33733] + MEM[33758];
assign MEM[41709] = MEM[33734] + MEM[33737];
assign MEM[41710] = MEM[33735] + MEM[33747];
assign MEM[41711] = MEM[33737] + MEM[33850];
assign MEM[41712] = MEM[33738] + MEM[33744];
assign MEM[41713] = MEM[33739] + MEM[33741];
assign MEM[41714] = MEM[33739] + MEM[33805];
assign MEM[41715] = MEM[33740] + MEM[33743];
assign MEM[41716] = MEM[33740] + MEM[33756];
assign MEM[41717] = MEM[33742] + MEM[33760];
assign MEM[41718] = MEM[33742] + MEM[33815];
assign MEM[41719] = MEM[33743] + MEM[33752];
assign MEM[41720] = MEM[33744] + MEM[33751];
assign MEM[41721] = MEM[33745] + MEM[33795];
assign MEM[41722] = MEM[33746] + MEM[33752];
assign MEM[41723] = MEM[33747] + MEM[33769];
assign MEM[41724] = MEM[33748] + MEM[33774];
assign MEM[41725] = MEM[33749] + MEM[33771];
assign MEM[41726] = MEM[33751] + MEM[33771];
assign MEM[41727] = MEM[33753] + MEM[33779];
assign MEM[41728] = MEM[33753] + MEM[33848];
assign MEM[41729] = MEM[33754] + MEM[33792];
assign MEM[41730] = MEM[33754] + MEM[33801];
assign MEM[41731] = MEM[33755] + MEM[33772];
assign MEM[41732] = MEM[33755] + MEM[33861];
assign MEM[41733] = MEM[33756] + MEM[33799];
assign MEM[41734] = MEM[33757] + MEM[33768];
assign MEM[41735] = MEM[33757] + MEM[33789];
assign MEM[41736] = MEM[33758] + MEM[33759];
assign MEM[41737] = MEM[33761] + MEM[33804];
assign MEM[41738] = MEM[33764] + MEM[33767];
assign MEM[41739] = MEM[33764] + MEM[33773];
assign MEM[41740] = MEM[33766] + MEM[33777];
assign MEM[41741] = MEM[33767] + MEM[33784];
assign MEM[41742] = MEM[33768] + MEM[33775];
assign MEM[41743] = MEM[33769] + MEM[33794];
assign MEM[41744] = MEM[33772] + MEM[33783];
assign MEM[41745] = MEM[33773] + MEM[33807];
assign MEM[41746] = MEM[33774] + MEM[33848];
assign MEM[41747] = MEM[33776] + MEM[33801];
assign MEM[41748] = MEM[33776] + MEM[33810];
assign MEM[41749] = MEM[33778] + MEM[33786];
assign MEM[41750] = MEM[33778] + MEM[33854];
assign MEM[41751] = MEM[33779] + MEM[33782];
assign MEM[41752] = MEM[33780] + MEM[33785];
assign MEM[41753] = MEM[33780] + MEM[33807];
assign MEM[41754] = MEM[33781] + MEM[33790];
assign MEM[41755] = MEM[33781] + MEM[33847];
assign MEM[41756] = MEM[33782] + MEM[33809];
assign MEM[41757] = MEM[33783] + MEM[33791];
assign MEM[41758] = MEM[33784] + MEM[33858];
assign MEM[41759] = MEM[33785] + MEM[33788];
assign MEM[41760] = MEM[33786] + MEM[33822];
assign MEM[41761] = MEM[33787] + MEM[33803];
assign MEM[41762] = MEM[33788] + MEM[33882];
assign MEM[41763] = MEM[33790] + MEM[33816];
assign MEM[41764] = MEM[33791] + MEM[33819];
assign MEM[41765] = MEM[33792] + MEM[33823];
assign MEM[41766] = MEM[33793] + MEM[33796];
assign MEM[41767] = MEM[33793] + MEM[33830];
assign MEM[41768] = MEM[33794] + MEM[33800];
assign MEM[41769] = MEM[33795] + MEM[33909];
assign MEM[41770] = MEM[33796] + MEM[33878];
assign MEM[41771] = MEM[33797] + MEM[33799];
assign MEM[41772] = MEM[33797] + MEM[33850];
assign MEM[41773] = MEM[33798] + MEM[33862];
assign MEM[41774] = MEM[33800] + MEM[33811];
assign MEM[41775] = MEM[33802] + MEM[33826];
assign MEM[41776] = MEM[33802] + MEM[33884];
assign MEM[41777] = MEM[33803] + MEM[33812];
assign MEM[41778] = MEM[33804] + MEM[33806];
assign MEM[41779] = MEM[33805] + MEM[33814];
assign MEM[41780] = MEM[33806] + MEM[33834];
assign MEM[41781] = MEM[33808] + MEM[33813];
assign MEM[41782] = MEM[33808] + MEM[33865];
assign MEM[41783] = MEM[33809] + MEM[33817];
assign MEM[41784] = MEM[33810] + MEM[33866];
assign MEM[41785] = MEM[33811] + MEM[33814];
assign MEM[41786] = MEM[33813] + MEM[33843];
assign MEM[41787] = MEM[33815] + MEM[33819];
assign MEM[41788] = MEM[33816] + MEM[33836];
assign MEM[41789] = MEM[33817] + MEM[33852];
assign MEM[41790] = MEM[33818] + MEM[33851];
assign MEM[41791] = MEM[33818] + MEM[33888];
assign MEM[41792] = MEM[33820] + MEM[33825];
assign MEM[41793] = MEM[33820] + MEM[33837];
assign MEM[41794] = MEM[33821] + MEM[33838];
assign MEM[41795] = MEM[33821] + MEM[33921];
assign MEM[41796] = MEM[33822] + MEM[33853];
assign MEM[41797] = MEM[33823] + MEM[33833];
assign MEM[41798] = MEM[33824] + MEM[33831];
assign MEM[41799] = MEM[33824] + MEM[33835];
assign MEM[41800] = MEM[33825] + MEM[33834];
assign MEM[41801] = MEM[33826] + MEM[33880];
assign MEM[41802] = MEM[33827] + MEM[33835];
assign MEM[41803] = MEM[33827] + MEM[33873];
assign MEM[41804] = MEM[33828] + MEM[33840];
assign MEM[41805] = MEM[33828] + MEM[33847];
assign MEM[41806] = MEM[33829] + MEM[33857];
assign MEM[41807] = MEM[33829] + MEM[33860];
assign MEM[41808] = MEM[33830] + MEM[33849];
assign MEM[41809] = MEM[33831] + MEM[33925];
assign MEM[41810] = MEM[33832] + MEM[33839];
assign MEM[41811] = MEM[33832] + MEM[33875];
assign MEM[41812] = MEM[33833] + MEM[33953];
assign MEM[41813] = MEM[33836] + MEM[33841];
assign MEM[41814] = MEM[33837] + MEM[33940];
assign MEM[41815] = MEM[33838] + MEM[33887];
assign MEM[41816] = MEM[33839] + MEM[33938];
assign MEM[41817] = MEM[33840] + MEM[33844];
assign MEM[41818] = MEM[33842] + MEM[33876];
assign MEM[41819] = MEM[33842] + MEM[33974];
assign MEM[41820] = MEM[33843] + MEM[33908];
assign MEM[41821] = MEM[33844] + MEM[33858];
assign MEM[41822] = MEM[33845] + MEM[33887];
assign MEM[41823] = MEM[33845] + MEM[33889];
assign MEM[41824] = MEM[33846] + MEM[33852];
assign MEM[41825] = MEM[33846] + MEM[33860];
assign MEM[41826] = MEM[33849] + MEM[33853];
assign MEM[41827] = MEM[33851] + MEM[33868];
assign MEM[41828] = MEM[33854] + MEM[33885];
assign MEM[41829] = MEM[33856] + MEM[33864];
assign MEM[41830] = MEM[33856] + MEM[33904];
assign MEM[41831] = MEM[33857] + MEM[33870];
assign MEM[41832] = MEM[33859] + MEM[33879];
assign MEM[41833] = MEM[33859] + MEM[33891];
assign MEM[41834] = MEM[33861] + MEM[33882];
assign MEM[41835] = MEM[33862] + MEM[34052];
assign MEM[41836] = MEM[33863] + MEM[33906];
assign MEM[41837] = MEM[33863] + MEM[33913];
assign MEM[41838] = MEM[33864] + MEM[33867];
assign MEM[41839] = MEM[33865] + MEM[33871];
assign MEM[41840] = MEM[33866] + MEM[33889];
assign MEM[41841] = MEM[33867] + MEM[33872];
assign MEM[41842] = MEM[33868] + MEM[33890];
assign MEM[41843] = MEM[33869] + MEM[33891];
assign MEM[41844] = MEM[33869] + MEM[33929];
assign MEM[41845] = MEM[33870] + MEM[33908];
assign MEM[41846] = MEM[33871] + MEM[33883];
assign MEM[41847] = MEM[33872] + MEM[33886];
assign MEM[41848] = MEM[33873] + MEM[33881];
assign MEM[41849] = MEM[33874] + MEM[33877];
assign MEM[41850] = MEM[33874] + MEM[33912];
assign MEM[41851] = MEM[33875] + MEM[33876];
assign MEM[41852] = MEM[33877] + MEM[33890];
assign MEM[41853] = MEM[33878] + MEM[33895];
assign MEM[41854] = MEM[33879] + MEM[33903];
assign MEM[41855] = MEM[33880] + MEM[33904];
assign MEM[41856] = MEM[33881] + MEM[33900];
assign MEM[41857] = MEM[33883] + MEM[33970];
assign MEM[41858] = MEM[33884] + MEM[33983];
assign MEM[41859] = MEM[33885] + MEM[33915];
assign MEM[41860] = MEM[33886] + MEM[33926];
assign MEM[41861] = MEM[33888] + MEM[33927];
assign MEM[41862] = MEM[33892] + MEM[33898];
assign MEM[41863] = MEM[33892] + MEM[33915];
assign MEM[41864] = MEM[33893] + MEM[33919];
assign MEM[41865] = MEM[33893] + MEM[33967];
assign MEM[41866] = MEM[33894] + MEM[33896];
assign MEM[41867] = MEM[33894] + MEM[33898];
assign MEM[41868] = MEM[33895] + MEM[33902];
assign MEM[41869] = MEM[33896] + MEM[33907];
assign MEM[41870] = MEM[33897] + MEM[33903];
assign MEM[41871] = MEM[33897] + MEM[33988];
assign MEM[41872] = MEM[33899] + MEM[33902];
assign MEM[41873] = MEM[33899] + MEM[33917];
assign MEM[41874] = MEM[33900] + MEM[33910];
assign MEM[41875] = MEM[33901] + MEM[33918];
assign MEM[41876] = MEM[33901] + MEM[33980];
assign MEM[41877] = MEM[33905] + MEM[33906];
assign MEM[41878] = MEM[33905] + MEM[33914];
assign MEM[41879] = MEM[33907] + MEM[33910];
assign MEM[41880] = MEM[33909] + MEM[33918];
assign MEM[41881] = MEM[33911] + MEM[33960];
assign MEM[41882] = MEM[33911] + MEM[34039];
assign MEM[41883] = MEM[33912] + MEM[33916];
assign MEM[41884] = MEM[33913] + MEM[34101];
assign MEM[41885] = MEM[33914] + MEM[33951];
assign MEM[41886] = MEM[33916] + MEM[33924];
assign MEM[41887] = MEM[33917] + MEM[33942];
assign MEM[41888] = MEM[33920] + MEM[33979];
assign MEM[41889] = MEM[33922] + MEM[34056];
assign MEM[41890] = MEM[33923] + MEM[33933];
assign MEM[41891] = MEM[33928] + MEM[34002];
assign MEM[41892] = MEM[33930] + MEM[33968];
assign MEM[41893] = MEM[33931] + MEM[34023];
assign MEM[41894] = MEM[33932] + MEM[34119];
assign MEM[41895] = MEM[33934] + MEM[33989];
assign MEM[41896] = MEM[33935] + MEM[34029];
assign MEM[41897] = MEM[33936] + MEM[34041];
assign MEM[41898] = MEM[33937] + MEM[33972];
assign MEM[41899] = MEM[33939] + MEM[34034];
assign MEM[41900] = MEM[33941] + MEM[34018];
assign MEM[41901] = MEM[33943] + MEM[33984];
assign MEM[41902] = MEM[33944] + MEM[34009];
assign MEM[41903] = MEM[33945] + MEM[34017];
assign MEM[41904] = MEM[33946] + MEM[34013];
assign MEM[41905] = MEM[33947] + MEM[34081];
assign MEM[41906] = MEM[33948] + MEM[34003];
assign MEM[41907] = MEM[33949] + MEM[33996];
assign MEM[41908] = MEM[33950] + MEM[34084];
assign MEM[41909] = MEM[33952] + MEM[34038];
assign MEM[41910] = MEM[33954] + MEM[34051];
assign MEM[41911] = MEM[33955] + MEM[34026];
assign MEM[41912] = MEM[33956] + MEM[34050];
assign MEM[41913] = MEM[33957] + MEM[33987];
assign MEM[41914] = MEM[33958] + MEM[34096];
assign MEM[41915] = MEM[33959] + MEM[34001];
assign MEM[41916] = MEM[33961] + MEM[34058];
assign MEM[41917] = MEM[33962] + MEM[34064];
assign MEM[41918] = MEM[33963] + MEM[34077];
assign MEM[41919] = MEM[33964] + MEM[34010];
assign MEM[41920] = MEM[33965] + MEM[34024];
assign MEM[41921] = MEM[33966] + MEM[33985];
assign MEM[41922] = MEM[33969] + MEM[33981];
assign MEM[41923] = MEM[33971] + MEM[34006];
assign MEM[41924] = MEM[33973] + MEM[34044];
assign MEM[41925] = MEM[33975] + MEM[33998];
assign MEM[41926] = MEM[33976] + MEM[34021];
assign MEM[41927] = MEM[33977] + MEM[34078];
assign MEM[41928] = MEM[33978] + MEM[34011];
assign MEM[41929] = MEM[33982] + MEM[34043];
assign MEM[41930] = MEM[33986] + MEM[34066];
assign MEM[41931] = MEM[33990] + MEM[34012];
assign MEM[41932] = MEM[33991] + MEM[34027];
assign MEM[41933] = MEM[33992] + MEM[34020];
assign MEM[41934] = MEM[33993] + MEM[34059];
assign MEM[41935] = MEM[33994] + MEM[33999];
assign MEM[41936] = MEM[33995] + MEM[34146];
assign MEM[41937] = MEM[33997] + MEM[34008];
assign MEM[41938] = MEM[34000] + MEM[34091];
assign MEM[41939] = MEM[34004] + MEM[34054];
assign MEM[41940] = MEM[34005] + MEM[34040];
assign MEM[41941] = MEM[34007] + MEM[34045];
assign MEM[41942] = MEM[34014] + MEM[34022];
assign MEM[41943] = MEM[34015] + MEM[34068];
assign MEM[41944] = MEM[34016] + MEM[34053];
assign MEM[41945] = MEM[34019] + MEM[34106];
assign MEM[41946] = MEM[34025] + MEM[34156];
assign MEM[41947] = MEM[34028] + MEM[34042];
assign MEM[41948] = MEM[34030] + MEM[34150];
assign MEM[41949] = MEM[34031] + MEM[34152];
assign MEM[41950] = MEM[34032] + MEM[34093];
assign MEM[41951] = MEM[34033] + MEM[34189];
assign MEM[41952] = MEM[34035] + MEM[34060];
assign MEM[41953] = MEM[34036] + MEM[34067];
assign MEM[41954] = MEM[34037] + MEM[34063];
assign MEM[41955] = MEM[34046] + MEM[34112];
assign MEM[41956] = MEM[34047] + MEM[34243];
assign MEM[41957] = MEM[34048] + MEM[34083];
assign MEM[41958] = MEM[34049] + MEM[34069];
assign MEM[41959] = MEM[34055] + MEM[34065];
assign MEM[41960] = MEM[34057] + MEM[34158];
assign MEM[41961] = MEM[34061] + MEM[34075];
assign MEM[41962] = MEM[34062] + MEM[34129];
assign MEM[41963] = MEM[34070] + MEM[34073];
assign MEM[41964] = MEM[34071] + MEM[34159];
assign MEM[41965] = MEM[34072] + MEM[34160];
assign MEM[41966] = MEM[34074] + MEM[34114];
assign MEM[41967] = MEM[34076] + MEM[34161];
assign MEM[41968] = MEM[34079] + MEM[34198];
assign MEM[41969] = MEM[34080] + MEM[34144];
assign MEM[41970] = MEM[34082] + MEM[34131];
assign MEM[41971] = MEM[34085] + MEM[34171];
assign MEM[41972] = MEM[34086] + MEM[34090];
assign MEM[41973] = MEM[34087] + MEM[34169];
assign MEM[41974] = MEM[34088] + MEM[34143];
assign MEM[41975] = MEM[34089] + MEM[34162];
assign MEM[41976] = MEM[34092] + MEM[34109];
assign MEM[41977] = MEM[34094] + MEM[34132];
assign MEM[41978] = MEM[34095] + MEM[34124];
assign MEM[41979] = MEM[34097] + MEM[34100];
assign MEM[41980] = MEM[34098] + MEM[34145];
assign MEM[41981] = MEM[34099] + MEM[34141];
assign MEM[41982] = MEM[34102] + MEM[34194];
assign MEM[41983] = MEM[34103] + MEM[34173];
assign MEM[41984] = MEM[34104] + MEM[34127];
assign MEM[41985] = MEM[34105] + MEM[34116];
assign MEM[41986] = MEM[34107] + MEM[34135];
assign MEM[41987] = MEM[34108] + MEM[34187];
assign MEM[41988] = MEM[34110] + MEM[34142];
assign MEM[41989] = MEM[34111] + MEM[34136];
assign MEM[41990] = MEM[34113] + MEM[34212];
assign MEM[41991] = MEM[34115] + MEM[34154];
assign MEM[41992] = MEM[34117] + MEM[34120];
assign MEM[41993] = MEM[34118] + MEM[34165];
assign MEM[41994] = MEM[34121] + MEM[34337];
assign MEM[41995] = MEM[34122] + MEM[34175];
assign MEM[41996] = MEM[34123] + MEM[34345];
assign MEM[41997] = MEM[34125] + MEM[34149];
assign MEM[41998] = MEM[34126] + MEM[34237];
assign MEM[41999] = MEM[34128] + MEM[34207];
assign MEM[42000] = MEM[34130] + MEM[34134];
assign MEM[42001] = MEM[34133] + MEM[34166];
assign MEM[42002] = MEM[34137] + MEM[34206];
assign MEM[42003] = MEM[34138] + MEM[34172];
assign MEM[42004] = MEM[34139] + MEM[34163];
assign MEM[42005] = MEM[34140] + MEM[34247];
assign MEM[42006] = MEM[34147] + MEM[34215];
assign MEM[42007] = MEM[34148] + MEM[34209];
assign MEM[42008] = MEM[34151] + MEM[34234];
assign MEM[42009] = MEM[34153] + MEM[34239];
assign MEM[42010] = MEM[34155] + MEM[34211];
assign MEM[42011] = MEM[34157] + MEM[34220];
assign MEM[42012] = MEM[34164] + MEM[34199];
assign MEM[42013] = MEM[34167] + MEM[34168];
assign MEM[42014] = MEM[34170] + MEM[34200];
assign MEM[42015] = MEM[34174] + MEM[34258];
assign MEM[42016] = MEM[34176] + MEM[34190];
assign MEM[42017] = MEM[34177] + MEM[34208];
assign MEM[42018] = MEM[34178] + MEM[34233];
assign MEM[42019] = MEM[34179] + MEM[34289];
assign MEM[42020] = MEM[34180] + MEM[34214];
assign MEM[42021] = MEM[34181] + MEM[34221];
assign MEM[42022] = MEM[34182] + MEM[34205];
assign MEM[42023] = MEM[34183] + MEM[34312];
assign MEM[42024] = MEM[34184] + MEM[34196];
assign MEM[42025] = MEM[34185] + MEM[34257];
assign MEM[42026] = MEM[34186] + MEM[34281];
assign MEM[42027] = MEM[34188] + MEM[34349];
assign MEM[42028] = MEM[34191] + MEM[34364];
assign MEM[42029] = MEM[34192] + MEM[34296];
assign MEM[42030] = MEM[34193] + MEM[34226];
assign MEM[42031] = MEM[34195] + MEM[34437];
assign MEM[42032] = MEM[34197] + MEM[34235];
assign MEM[42033] = MEM[34201] + MEM[34429];
assign MEM[42034] = MEM[34202] + MEM[34231];
assign MEM[42035] = MEM[34203] + MEM[34260];
assign MEM[42036] = MEM[34204] + MEM[34236];
assign MEM[42037] = MEM[34210] + MEM[34300];
assign MEM[42038] = MEM[34213] + MEM[34240];
assign MEM[42039] = MEM[34216] + MEM[34261];
assign MEM[42040] = MEM[34217] + MEM[34264];
assign MEM[42041] = MEM[34218] + MEM[34330];
assign MEM[42042] = MEM[34219] + MEM[34263];
assign MEM[42043] = MEM[34222] + MEM[34254];
assign MEM[42044] = MEM[34223] + MEM[34250];
assign MEM[42045] = MEM[34224] + MEM[34302];
assign MEM[42046] = MEM[34225] + MEM[34321];
assign MEM[42047] = MEM[34227] + MEM[34417];
assign MEM[42048] = MEM[34228] + MEM[34266];
assign MEM[42049] = MEM[34229] + MEM[34310];
assign MEM[42050] = MEM[34230] + MEM[34241];
assign MEM[42051] = MEM[34232] + MEM[34354];
assign MEM[42052] = MEM[34238] + MEM[34291];
assign MEM[42053] = MEM[34242] + MEM[34313];
assign MEM[42054] = MEM[34244] + MEM[34249];
assign MEM[42055] = MEM[34245] + MEM[34332];
assign MEM[42056] = MEM[34246] + MEM[34316];
assign MEM[42057] = MEM[34248] + MEM[34294];
assign MEM[42058] = MEM[34251] + MEM[34369];
assign MEM[42059] = MEM[34252] + MEM[34297];
assign MEM[42060] = MEM[34253] + MEM[34352];
assign MEM[42061] = MEM[34255] + MEM[34267];
assign MEM[42062] = MEM[34256] + MEM[34287];
assign MEM[42063] = MEM[34259] + MEM[34329];
assign MEM[42064] = MEM[34262] + MEM[34315];
assign MEM[42065] = MEM[34265] + MEM[34326];
assign MEM[42066] = MEM[34268] + MEM[34280];
assign MEM[42067] = MEM[34269] + MEM[34301];
assign MEM[42068] = MEM[34270] + MEM[34308];
assign MEM[42069] = MEM[34271] + MEM[34277];
assign MEM[42070] = MEM[34272] + MEM[34305];
assign MEM[42071] = MEM[34273] + MEM[34397];
assign MEM[42072] = MEM[34274] + MEM[34311];
assign MEM[42073] = MEM[34275] + MEM[34357];
assign MEM[42074] = MEM[34276] + MEM[34338];
assign MEM[42075] = MEM[34278] + MEM[34314];
assign MEM[42076] = MEM[34279] + MEM[34318];
assign MEM[42077] = MEM[34282] + MEM[34320];
assign MEM[42078] = MEM[34283] + MEM[34356];
assign MEM[42079] = MEM[34284] + MEM[34390];
assign MEM[42080] = MEM[34285] + MEM[34394];
assign MEM[42081] = MEM[34286] + MEM[34453];
assign MEM[42082] = MEM[34288] + MEM[34420];
assign MEM[42083] = MEM[34290] + MEM[34292];
assign MEM[42084] = MEM[34293] + MEM[34307];
assign MEM[42085] = MEM[34295] + MEM[34327];
assign MEM[42086] = MEM[34298] + MEM[34463];
assign MEM[42087] = MEM[34299] + MEM[34387];
assign MEM[42088] = MEM[34303] + MEM[34335];
assign MEM[42089] = MEM[34304] + MEM[34348];
assign MEM[42090] = MEM[34306] + MEM[34392];
assign MEM[42091] = MEM[34309] + MEM[34346];
assign MEM[42092] = MEM[34317] + MEM[34374];
assign MEM[42093] = MEM[34319] + MEM[34336];
assign MEM[42094] = MEM[34322] + MEM[34358];
assign MEM[42095] = MEM[34323] + MEM[34373];
assign MEM[42096] = MEM[34324] + MEM[34341];
assign MEM[42097] = MEM[34325] + MEM[34432];
assign MEM[42098] = MEM[34328] + MEM[34343];
assign MEM[42099] = MEM[34331] + MEM[34351];
assign MEM[42100] = MEM[34333] + MEM[34359];
assign MEM[42101] = MEM[34334] + MEM[34376];
assign MEM[42102] = MEM[34339] + MEM[34382];
assign MEM[42103] = MEM[34340] + MEM[34347];
assign MEM[42104] = MEM[34342] + MEM[34413];
assign MEM[42105] = MEM[34344] + MEM[34370];
assign MEM[42106] = MEM[34350] + MEM[34405];
assign MEM[42107] = MEM[34353] + MEM[34408];
assign MEM[42108] = MEM[34355] + MEM[34419];
assign MEM[42109] = MEM[34360] + MEM[34368];
assign MEM[42110] = MEM[34361] + MEM[34388];
assign MEM[42111] = MEM[34362] + MEM[34385];
assign MEM[42112] = MEM[34363] + MEM[34502];
assign MEM[42113] = MEM[34365] + MEM[34399];
assign MEM[42114] = MEM[34366] + MEM[34367];
assign MEM[42115] = MEM[34371] + MEM[34468];
assign MEM[42116] = MEM[34372] + MEM[34427];
assign MEM[42117] = MEM[34375] + MEM[34396];
assign MEM[42118] = MEM[34377] + MEM[34411];
assign MEM[42119] = MEM[34378] + MEM[34416];
assign MEM[42120] = MEM[34379] + MEM[34464];
assign MEM[42121] = MEM[34380] + MEM[34527];
assign MEM[42122] = MEM[34381] + MEM[34401];
assign MEM[42123] = MEM[34383] + MEM[34421];
assign MEM[42124] = MEM[34384] + MEM[34491];
assign MEM[42125] = MEM[34386] + MEM[34454];
assign MEM[42126] = MEM[34389] + MEM[34403];
assign MEM[42127] = MEM[34391] + MEM[34410];
assign MEM[42128] = MEM[34393] + MEM[34439];
assign MEM[42129] = MEM[34395] + MEM[34412];
assign MEM[42130] = MEM[34398] + MEM[34406];
assign MEM[42131] = MEM[34400] + MEM[34436];
assign MEM[42132] = MEM[34402] + MEM[34449];
assign MEM[42133] = MEM[34404] + MEM[34474];
assign MEM[42134] = MEM[34407] + MEM[34554];
assign MEM[42135] = MEM[34409] + MEM[34448];
assign MEM[42136] = MEM[34414] + MEM[34441];
assign MEM[42137] = MEM[34415] + MEM[34455];
assign MEM[42138] = MEM[34418] + MEM[34484];
assign MEM[42139] = MEM[34422] + MEM[34533];
assign MEM[42140] = MEM[34423] + MEM[34529];
assign MEM[42141] = MEM[34424] + MEM[34466];
assign MEM[42142] = MEM[34425] + MEM[34447];
assign MEM[42143] = MEM[34426] + MEM[34445];
assign MEM[42144] = MEM[34428] + MEM[34539];
assign MEM[42145] = MEM[34430] + MEM[34510];
assign MEM[42146] = MEM[34431] + MEM[34440];
assign MEM[42147] = MEM[34433] + MEM[34496];
assign MEM[42148] = MEM[34434] + MEM[34472];
assign MEM[42149] = MEM[34435] + MEM[34481];
assign MEM[42150] = MEM[34438] + MEM[34475];
assign MEM[42151] = MEM[34442] + MEM[34458];
assign MEM[42152] = MEM[34443] + MEM[34519];
assign MEM[42153] = MEM[34444] + MEM[34495];
assign MEM[42154] = MEM[34446] + MEM[34633];
assign MEM[42155] = MEM[34450] + MEM[34461];
assign MEM[42156] = MEM[34451] + MEM[34561];
assign MEM[42157] = MEM[34452] + MEM[34482];
assign MEM[42158] = MEM[34456] + MEM[34579];
assign MEM[42159] = MEM[34457] + MEM[34479];
assign MEM[42160] = MEM[34459] + MEM[34476];
assign MEM[42161] = MEM[34460] + MEM[34511];
assign MEM[42162] = MEM[34462] + MEM[34516];
assign MEM[42163] = MEM[34465] + MEM[34509];
assign MEM[42164] = MEM[34467] + MEM[34505];
assign MEM[42165] = MEM[34469] + MEM[34512];
assign MEM[42166] = MEM[34470] + MEM[34487];
assign MEM[42167] = MEM[34471] + MEM[34528];
assign MEM[42168] = MEM[34473] + MEM[34480];
assign MEM[42169] = MEM[34477] + MEM[34540];
assign MEM[42170] = MEM[34478] + MEM[34553];
assign MEM[42171] = MEM[34483] + MEM[34611];
assign MEM[42172] = MEM[34485] + MEM[34549];
assign MEM[42173] = MEM[34486] + MEM[34585];
assign MEM[42174] = MEM[34488] + MEM[34701];
assign MEM[42175] = MEM[34489] + MEM[34518];
assign MEM[42176] = MEM[34490] + MEM[34501];
assign MEM[42177] = MEM[34492] + MEM[34504];
assign MEM[42178] = MEM[34493] + MEM[34559];
assign MEM[42179] = MEM[34494] + MEM[34541];
assign MEM[42180] = MEM[34497] + MEM[34506];
assign MEM[42181] = MEM[34498] + MEM[34551];
assign MEM[42182] = MEM[34499] + MEM[34530];
assign MEM[42183] = MEM[34500] + MEM[34576];
assign MEM[42184] = MEM[34503] + MEM[34524];
assign MEM[42185] = MEM[34507] + MEM[34629];
assign MEM[42186] = MEM[34508] + MEM[34534];
assign MEM[42187] = MEM[34513] + MEM[34622];
assign MEM[42188] = MEM[34514] + MEM[34597];
assign MEM[42189] = MEM[34515] + MEM[34584];
assign MEM[42190] = MEM[34517] + MEM[34543];
assign MEM[42191] = MEM[34520] + MEM[34535];
assign MEM[42192] = MEM[34521] + MEM[34625];
assign MEM[42193] = MEM[34522] + MEM[34548];
assign MEM[42194] = MEM[34523] + MEM[34580];
assign MEM[42195] = MEM[34525] + MEM[34569];
assign MEM[42196] = MEM[34526] + MEM[34562];
assign MEM[42197] = MEM[34531] + MEM[34555];
assign MEM[42198] = MEM[34532] + MEM[34616];
assign MEM[42199] = MEM[34536] + MEM[34538];
assign MEM[42200] = MEM[34537] + MEM[34610];
assign MEM[42201] = MEM[34542] + MEM[34608];
assign MEM[42202] = MEM[34544] + MEM[34696];
assign MEM[42203] = MEM[34545] + MEM[34617];
assign MEM[42204] = MEM[34546] + MEM[34592];
assign MEM[42205] = MEM[34547] + MEM[34729];
assign MEM[42206] = MEM[34550] + MEM[34602];
assign MEM[42207] = MEM[34552] + MEM[34577];
assign MEM[42208] = MEM[34556] + MEM[34609];
assign MEM[42209] = MEM[34557] + MEM[34598];
assign MEM[42210] = MEM[34558] + MEM[34634];
assign MEM[42211] = MEM[34560] + MEM[34568];
assign MEM[42212] = MEM[34563] + MEM[34620];
assign MEM[42213] = MEM[34564] + MEM[34578];
assign MEM[42214] = MEM[34565] + MEM[34626];
assign MEM[42215] = MEM[34566] + MEM[34640];
assign MEM[42216] = MEM[34567] + MEM[34657];
assign MEM[42217] = MEM[34570] + MEM[34644];
assign MEM[42218] = MEM[34571] + MEM[34720];
assign MEM[42219] = MEM[34572] + MEM[34581];
assign MEM[42220] = MEM[34573] + MEM[34661];
assign MEM[42221] = MEM[34574] + MEM[34646];
assign MEM[42222] = MEM[34575] + MEM[34824];
assign MEM[42223] = MEM[34582] + MEM[34651];
assign MEM[42224] = MEM[34583] + MEM[34655];
assign MEM[42225] = MEM[34586] + MEM[34702];
assign MEM[42226] = MEM[34587] + MEM[34638];
assign MEM[42227] = MEM[34588] + MEM[34596];
assign MEM[42228] = MEM[34589] + MEM[34645];
assign MEM[42229] = MEM[34590] + MEM[34636];
assign MEM[42230] = MEM[34591] + MEM[34664];
assign MEM[42231] = MEM[34593] + MEM[34603];
assign MEM[42232] = MEM[34594] + MEM[34612];
assign MEM[42233] = MEM[34595] + MEM[34606];
assign MEM[42234] = MEM[34599] + MEM[34641];
assign MEM[42235] = MEM[34600] + MEM[34614];
assign MEM[42236] = MEM[34601] + MEM[34709];
assign MEM[42237] = MEM[34604] + MEM[34619];
assign MEM[42238] = MEM[34605] + MEM[34628];
assign MEM[42239] = MEM[34607] + MEM[34668];
assign MEM[42240] = MEM[34613] + MEM[34690];
assign MEM[42241] = MEM[34615] + MEM[34707];
assign MEM[42242] = MEM[34618] + MEM[34687];
assign MEM[42243] = MEM[34621] + MEM[34624];
assign MEM[42244] = MEM[34623] + MEM[34695];
assign MEM[42245] = MEM[34627] + MEM[34773];
assign MEM[42246] = MEM[34630] + MEM[34708];
assign MEM[42247] = MEM[34631] + MEM[34671];
assign MEM[42248] = MEM[34632] + MEM[34694];
assign MEM[42249] = MEM[34635] + MEM[34648];
assign MEM[42250] = MEM[34637] + MEM[34643];
assign MEM[42251] = MEM[34639] + MEM[34725];
assign MEM[42252] = MEM[34642] + MEM[34742];
assign MEM[42253] = MEM[34647] + MEM[34705];
assign MEM[42254] = MEM[34649] + MEM[34670];
assign MEM[42255] = MEM[34650] + MEM[34684];
assign MEM[42256] = MEM[34652] + MEM[34697];
assign MEM[42257] = MEM[34653] + MEM[34706];
assign MEM[42258] = MEM[34654] + MEM[34746];
assign MEM[42259] = MEM[34656] + MEM[34672];
assign MEM[42260] = MEM[34658] + MEM[34737];
assign MEM[42261] = MEM[34659] + MEM[34804];
assign MEM[42262] = MEM[34660] + MEM[34692];
assign MEM[42263] = MEM[34662] + MEM[34731];
assign MEM[42264] = MEM[34663] + MEM[34734];
assign MEM[42265] = MEM[34665] + MEM[34712];
assign MEM[42266] = MEM[34666] + MEM[34673];
assign MEM[42267] = MEM[34667] + MEM[34783];
assign MEM[42268] = MEM[34669] + MEM[34739];
assign MEM[42269] = MEM[34674] + MEM[34747];
assign MEM[42270] = MEM[34675] + MEM[34721];
assign MEM[42271] = MEM[34676] + MEM[34727];
assign MEM[42272] = MEM[34677] + MEM[34719];
assign MEM[42273] = MEM[34678] + MEM[34780];
assign MEM[42274] = MEM[34679] + MEM[34843];
assign MEM[42275] = MEM[34680] + MEM[34724];
assign MEM[42276] = MEM[34681] + MEM[34726];
assign MEM[42277] = MEM[34682] + MEM[34704];
assign MEM[42278] = MEM[34683] + MEM[34743];
assign MEM[42279] = MEM[34685] + MEM[34749];
assign MEM[42280] = MEM[34686] + MEM[34900];
assign MEM[42281] = MEM[34688] + MEM[34777];
assign MEM[42282] = MEM[34689] + MEM[34738];
assign MEM[42283] = MEM[34691] + MEM[34764];
assign MEM[42284] = MEM[34693] + MEM[34840];
assign MEM[42285] = MEM[34698] + MEM[34735];
assign MEM[42286] = MEM[34699] + MEM[34771];
assign MEM[42287] = MEM[34700] + MEM[34748];
assign MEM[42288] = MEM[34703] + MEM[34789];
assign MEM[42289] = MEM[34710] + MEM[34753];
assign MEM[42290] = MEM[34711] + MEM[34745];
assign MEM[42291] = MEM[34713] + MEM[34766];
assign MEM[42292] = MEM[34714] + MEM[34740];
assign MEM[42293] = MEM[34715] + MEM[34756];
assign MEM[42294] = MEM[34716] + MEM[34723];
assign MEM[42295] = MEM[34717] + MEM[34794];
assign MEM[42296] = MEM[34718] + MEM[34758];
assign MEM[42297] = MEM[34722] + MEM[34761];
assign MEM[42298] = MEM[34728] + MEM[34744];
assign MEM[42299] = MEM[34730] + MEM[34852];
assign MEM[42300] = MEM[34732] + MEM[34925];
assign MEM[42301] = MEM[34733] + MEM[34938];
assign MEM[42302] = MEM[34736] + MEM[34838];
assign MEM[42303] = MEM[34741] + MEM[35051];
assign MEM[42304] = MEM[34750] + MEM[34793];
assign MEM[42305] = MEM[34751] + MEM[34796];
assign MEM[42306] = MEM[34752] + MEM[34814];
assign MEM[42307] = MEM[34754] + MEM[34782];
assign MEM[42308] = MEM[34755] + MEM[34781];
assign MEM[42309] = MEM[34757] + MEM[34832];
assign MEM[42310] = MEM[34759] + MEM[34774];
assign MEM[42311] = MEM[34760] + MEM[34821];
assign MEM[42312] = MEM[34762] + MEM[34842];
assign MEM[42313] = MEM[34763] + MEM[34950];
assign MEM[42314] = MEM[34765] + MEM[34788];
assign MEM[42315] = MEM[34767] + MEM[34792];
assign MEM[42316] = MEM[34768] + MEM[34785];
assign MEM[42317] = MEM[34769] + MEM[34811];
assign MEM[42318] = MEM[34770] + MEM[34901];
assign MEM[42319] = MEM[34772] + MEM[34815];
assign MEM[42320] = MEM[34775] + MEM[34798];
assign MEM[42321] = MEM[34776] + MEM[34826];
assign MEM[42322] = MEM[34778] + MEM[34904];
assign MEM[42323] = MEM[34779] + MEM[34819];
assign MEM[42324] = MEM[34784] + MEM[34846];
assign MEM[42325] = MEM[34786] + MEM[34791];
assign MEM[42326] = MEM[34787] + MEM[34825];
assign MEM[42327] = MEM[34790] + MEM[34841];
assign MEM[42328] = MEM[34795] + MEM[34837];
assign MEM[42329] = MEM[34797] + MEM[34834];
assign MEM[42330] = MEM[34799] + MEM[34885];
assign MEM[42331] = MEM[34800] + MEM[34907];
assign MEM[42332] = MEM[34801] + MEM[34827];
assign MEM[42333] = MEM[34802] + MEM[34816];
assign MEM[42334] = MEM[34803] + MEM[34855];
assign MEM[42335] = MEM[34805] + MEM[34856];
assign MEM[42336] = MEM[34806] + MEM[34829];
assign MEM[42337] = MEM[34807] + MEM[34929];
assign MEM[42338] = MEM[34808] + MEM[34857];
assign MEM[42339] = MEM[34809] + MEM[34899];
assign MEM[42340] = MEM[34810] + MEM[34873];
assign MEM[42341] = MEM[34812] + MEM[34866];
assign MEM[42342] = MEM[34813] + MEM[34920];
assign MEM[42343] = MEM[34817] + MEM[34862];
assign MEM[42344] = MEM[34818] + MEM[34930];
assign MEM[42345] = MEM[34820] + MEM[34891];
assign MEM[42346] = MEM[34822] + MEM[34871];
assign MEM[42347] = MEM[34823] + MEM[34882];
assign MEM[42348] = MEM[34828] + MEM[34897];
assign MEM[42349] = MEM[34830] + MEM[34909];
assign MEM[42350] = MEM[34831] + MEM[34916];
assign MEM[42351] = MEM[34833] + MEM[34848];
assign MEM[42352] = MEM[34835] + MEM[34968];
assign MEM[42353] = MEM[34836] + MEM[34884];
assign MEM[42354] = MEM[34839] + MEM[34875];
assign MEM[42355] = MEM[34844] + MEM[34989];
assign MEM[42356] = MEM[34845] + MEM[34880];
assign MEM[42357] = MEM[34847] + MEM[34887];
assign MEM[42358] = MEM[34849] + MEM[34854];
assign MEM[42359] = MEM[34850] + MEM[34924];
assign MEM[42360] = MEM[34851] + MEM[34954];
assign MEM[42361] = MEM[34853] + MEM[34869];
assign MEM[42362] = MEM[34858] + MEM[34898];
assign MEM[42363] = MEM[34859] + MEM[34926];
assign MEM[42364] = MEM[34860] + MEM[34889];
assign MEM[42365] = MEM[34861] + MEM[34985];
assign MEM[42366] = MEM[34863] + MEM[34910];
assign MEM[42367] = MEM[34864] + MEM[34908];
assign MEM[42368] = MEM[34865] + MEM[34918];
assign MEM[42369] = MEM[34867] + MEM[34883];
assign MEM[42370] = MEM[34868] + MEM[34942];
assign MEM[42371] = MEM[34870] + MEM[34905];
assign MEM[42372] = MEM[34872] + MEM[34964];
assign MEM[42373] = MEM[34874] + MEM[34876];
assign MEM[42374] = MEM[34877] + MEM[34911];
assign MEM[42375] = MEM[34878] + MEM[34959];
assign MEM[42376] = MEM[34879] + MEM[34935];
assign MEM[42377] = MEM[34881] + MEM[34982];
assign MEM[42378] = MEM[34886] + MEM[34917];
assign MEM[42379] = MEM[34888] + MEM[34979];
assign MEM[42380] = MEM[34890] + MEM[35111];
assign MEM[42381] = MEM[34892] + MEM[34983];
assign MEM[42382] = MEM[34893] + MEM[35005];
assign MEM[42383] = MEM[34894] + MEM[34956];
assign MEM[42384] = MEM[34895] + MEM[34945];
assign MEM[42385] = MEM[34896] + MEM[34977];
assign MEM[42386] = MEM[34902] + MEM[34963];
assign MEM[42387] = MEM[34903] + MEM[34914];
assign MEM[42388] = MEM[34906] + MEM[34915];
assign MEM[42389] = MEM[34912] + MEM[34941];
assign MEM[42390] = MEM[34913] + MEM[34934];
assign MEM[42391] = MEM[34919] + MEM[34984];
assign MEM[42392] = MEM[34921] + MEM[35113];
assign MEM[42393] = MEM[34922] + MEM[34932];
assign MEM[42394] = MEM[34923] + MEM[34990];
assign MEM[42395] = MEM[34927] + MEM[35074];
assign MEM[42396] = MEM[34928] + MEM[35058];
assign MEM[42397] = MEM[34931] + MEM[34969];
assign MEM[42398] = MEM[34933] + MEM[35000];
assign MEM[42399] = MEM[34936] + MEM[34999];
assign MEM[42400] = MEM[34937] + MEM[34978];
assign MEM[42401] = MEM[34939] + MEM[35039];
assign MEM[42402] = MEM[34940] + MEM[34976];
assign MEM[42403] = MEM[34943] + MEM[35013];
assign MEM[42404] = MEM[34944] + MEM[35015];
assign MEM[42405] = MEM[34946] + MEM[34998];
assign MEM[42406] = MEM[34947] + MEM[35023];
assign MEM[42407] = MEM[34948] + MEM[34970];
assign MEM[42408] = MEM[34949] + MEM[35012];
assign MEM[42409] = MEM[34951] + MEM[34972];
assign MEM[42410] = MEM[34952] + MEM[35029];
assign MEM[42411] = MEM[34953] + MEM[34960];
assign MEM[42412] = MEM[34955] + MEM[35034];
assign MEM[42413] = MEM[34957] + MEM[35032];
assign MEM[42414] = MEM[34958] + MEM[34988];
assign MEM[42415] = MEM[34961] + MEM[35108];
assign MEM[42416] = MEM[34962] + MEM[34986];
assign MEM[42417] = MEM[34965] + MEM[34997];
assign MEM[42418] = MEM[34966] + MEM[35024];
assign MEM[42419] = MEM[34967] + MEM[35060];
assign MEM[42420] = MEM[34971] + MEM[35036];
assign MEM[42421] = MEM[34973] + MEM[35188];
assign MEM[42422] = MEM[34974] + MEM[35002];
assign MEM[42423] = MEM[34975] + MEM[35094];
assign MEM[42424] = MEM[34980] + MEM[35044];
assign MEM[42425] = MEM[34981] + MEM[35091];
assign MEM[42426] = MEM[34987] + MEM[35089];
assign MEM[42427] = MEM[34991] + MEM[35010];
assign MEM[42428] = MEM[34992] + MEM[35014];
assign MEM[42429] = MEM[34993] + MEM[35028];
assign MEM[42430] = MEM[34994] + MEM[35020];
assign MEM[42431] = MEM[34995] + MEM[35030];
assign MEM[42432] = MEM[34996] + MEM[35031];
assign MEM[42433] = MEM[35001] + MEM[35123];
assign MEM[42434] = MEM[35003] + MEM[35017];
assign MEM[42435] = MEM[35004] + MEM[35008];
assign MEM[42436] = MEM[35006] + MEM[35079];
assign MEM[42437] = MEM[35007] + MEM[35083];
assign MEM[42438] = MEM[35009] + MEM[35056];
assign MEM[42439] = MEM[35011] + MEM[35057];
assign MEM[42440] = MEM[35016] + MEM[35112];
assign MEM[42441] = MEM[35018] + MEM[35053];
assign MEM[42442] = MEM[35019] + MEM[35037];
assign MEM[42443] = MEM[35021] + MEM[35070];
assign MEM[42444] = MEM[35022] + MEM[35049];
assign MEM[42445] = MEM[35025] + MEM[35282];
assign MEM[42446] = MEM[35026] + MEM[35084];
assign MEM[42447] = MEM[35027] + MEM[35077];
assign MEM[42448] = MEM[35033] + MEM[35048];
assign MEM[42449] = MEM[35035] + MEM[35090];
assign MEM[42450] = MEM[35038] + MEM[35142];
assign MEM[42451] = MEM[35040] + MEM[35180];
assign MEM[42452] = MEM[35041] + MEM[35129];
assign MEM[42453] = MEM[35042] + MEM[35069];
assign MEM[42454] = MEM[35043] + MEM[35149];
assign MEM[42455] = MEM[35045] + MEM[35055];
assign MEM[42456] = MEM[35046] + MEM[35216];
assign MEM[42457] = MEM[35047] + MEM[35078];
assign MEM[42458] = MEM[35050] + MEM[35109];
assign MEM[42459] = MEM[35052] + MEM[35076];
assign MEM[42460] = MEM[35054] + MEM[35101];
assign MEM[42461] = MEM[35059] + MEM[35116];
assign MEM[42462] = MEM[35061] + MEM[35140];
assign MEM[42463] = MEM[35062] + MEM[35175];
assign MEM[42464] = MEM[35063] + MEM[35066];
assign MEM[42465] = MEM[35064] + MEM[35088];
assign MEM[42466] = MEM[35065] + MEM[35086];
assign MEM[42467] = MEM[35067] + MEM[35117];
assign MEM[42468] = MEM[35068] + MEM[35127];
assign MEM[42469] = MEM[35071] + MEM[35155];
assign MEM[42470] = MEM[35072] + MEM[35183];
assign MEM[42471] = MEM[35073] + MEM[35143];
assign MEM[42472] = MEM[35075] + MEM[35095];
assign MEM[42473] = MEM[35080] + MEM[35102];
assign MEM[42474] = MEM[35081] + MEM[35119];
assign MEM[42475] = MEM[35082] + MEM[35097];
assign MEM[42476] = MEM[35085] + MEM[35310];
assign MEM[42477] = MEM[35087] + MEM[35159];
assign MEM[42478] = MEM[35092] + MEM[35106];
assign MEM[42479] = MEM[35093] + MEM[35137];
assign MEM[42480] = MEM[35096] + MEM[35191];
assign MEM[42481] = MEM[35098] + MEM[35195];
assign MEM[42482] = MEM[35099] + MEM[35125];
assign MEM[42483] = MEM[35100] + MEM[35165];
assign MEM[42484] = MEM[35103] + MEM[35139];
assign MEM[42485] = MEM[35104] + MEM[35174];
assign MEM[42486] = MEM[35105] + MEM[35151];
assign MEM[42487] = MEM[35107] + MEM[35264];
assign MEM[42488] = MEM[35110] + MEM[35168];
assign MEM[42489] = MEM[35114] + MEM[35152];
assign MEM[42490] = MEM[35115] + MEM[35164];
assign MEM[42491] = MEM[35118] + MEM[35171];
assign MEM[42492] = MEM[35120] + MEM[35178];
assign MEM[42493] = MEM[35121] + MEM[35187];
assign MEM[42494] = MEM[35122] + MEM[35157];
assign MEM[42495] = MEM[35124] + MEM[35287];
assign MEM[42496] = MEM[35126] + MEM[35141];
assign MEM[42497] = MEM[35128] + MEM[35312];
assign MEM[42498] = MEM[35130] + MEM[35240];
assign MEM[42499] = MEM[35131] + MEM[35213];
assign MEM[42500] = MEM[35132] + MEM[35177];
assign MEM[42501] = MEM[35133] + MEM[35212];
assign MEM[42502] = MEM[35134] + MEM[35146];
assign MEM[42503] = MEM[35135] + MEM[35307];
assign MEM[42504] = MEM[35136] + MEM[35145];
assign MEM[42505] = MEM[35138] + MEM[35182];
assign MEM[42506] = MEM[35144] + MEM[35203];
assign MEM[42507] = MEM[35147] + MEM[35179];
assign MEM[42508] = MEM[35148] + MEM[35205];
assign MEM[42509] = MEM[35150] + MEM[35245];
assign MEM[42510] = MEM[35153] + MEM[35356];
assign MEM[42511] = MEM[35154] + MEM[35207];
assign MEM[42512] = MEM[35156] + MEM[35252];
assign MEM[42513] = MEM[35158] + MEM[35272];
assign MEM[42514] = MEM[35160] + MEM[35176];
assign MEM[42515] = MEM[35161] + MEM[35221];
assign MEM[42516] = MEM[35162] + MEM[35173];
assign MEM[42517] = MEM[35163] + MEM[35199];
assign MEM[42518] = MEM[35166] + MEM[35228];
assign MEM[42519] = MEM[35167] + MEM[35342];
assign MEM[42520] = MEM[35169] + MEM[35241];
assign MEM[42521] = MEM[35170] + MEM[35248];
assign MEM[42522] = MEM[35172] + MEM[35194];
assign MEM[42523] = MEM[35181] + MEM[35277];
assign MEM[42524] = MEM[35184] + MEM[35292];
assign MEM[42525] = MEM[35185] + MEM[35209];
assign MEM[42526] = MEM[35186] + MEM[35247];
assign MEM[42527] = MEM[35189] + MEM[35267];
assign MEM[42528] = MEM[35190] + MEM[35284];
assign MEM[42529] = MEM[35192] + MEM[35255];
assign MEM[42530] = MEM[35193] + MEM[35269];
assign MEM[42531] = MEM[35196] + MEM[35233];
assign MEM[42532] = MEM[35197] + MEM[35332];
assign MEM[42533] = MEM[35198] + MEM[35211];
assign MEM[42534] = MEM[35200] + MEM[35259];
assign MEM[42535] = MEM[35201] + MEM[35275];
assign MEM[42536] = MEM[35202] + MEM[35242];
assign MEM[42537] = MEM[35204] + MEM[35273];
assign MEM[42538] = MEM[35206] + MEM[35218];
assign MEM[42539] = MEM[35208] + MEM[35263];
assign MEM[42540] = MEM[35210] + MEM[35230];
assign MEM[42541] = MEM[35214] + MEM[35229];
assign MEM[42542] = MEM[35215] + MEM[35232];
assign MEM[42543] = MEM[35217] + MEM[35250];
assign MEM[42544] = MEM[35219] + MEM[35262];
assign MEM[42545] = MEM[35220] + MEM[35234];
assign MEM[42546] = MEM[35222] + MEM[35305];
assign MEM[42547] = MEM[35223] + MEM[35261];
assign MEM[42548] = MEM[35224] + MEM[35349];
assign MEM[42549] = MEM[35225] + MEM[35283];
assign MEM[42550] = MEM[35226] + MEM[35260];
assign MEM[42551] = MEM[35227] + MEM[35246];
assign MEM[42552] = MEM[35231] + MEM[35296];
assign MEM[42553] = MEM[35235] + MEM[35270];
assign MEM[42554] = MEM[35236] + MEM[35289];
assign MEM[42555] = MEM[35237] + MEM[35291];
assign MEM[42556] = MEM[35238] + MEM[35357];
assign MEM[42557] = MEM[35239] + MEM[35300];
assign MEM[42558] = MEM[35243] + MEM[35367];
assign MEM[42559] = MEM[35244] + MEM[35352];
assign MEM[42560] = MEM[35249] + MEM[35323];
assign MEM[42561] = MEM[35251] + MEM[35359];
assign MEM[42562] = MEM[35253] + MEM[35453];
assign MEM[42563] = MEM[35254] + MEM[35302];
assign MEM[42564] = MEM[35256] + MEM[35304];
assign MEM[42565] = MEM[35257] + MEM[35274];
assign MEM[42566] = MEM[35258] + MEM[35322];
assign MEM[42567] = MEM[35265] + MEM[35343];
assign MEM[42568] = MEM[35266] + MEM[35466];
assign MEM[42569] = MEM[35268] + MEM[35407];
assign MEM[42570] = MEM[35271] + MEM[35317];
assign MEM[42571] = MEM[35276] + MEM[35301];
assign MEM[42572] = MEM[35278] + MEM[35386];
assign MEM[42573] = MEM[35279] + MEM[35358];
assign MEM[42574] = MEM[35280] + MEM[35330];
assign MEM[42575] = MEM[35281] + MEM[35295];
assign MEM[42576] = MEM[35285] + MEM[35346];
assign MEM[42577] = MEM[35286] + MEM[35294];
assign MEM[42578] = MEM[35288] + MEM[35396];
assign MEM[42579] = MEM[35290] + MEM[35320];
assign MEM[42580] = MEM[35293] + MEM[35309];
assign MEM[42581] = MEM[35297] + MEM[35347];
assign MEM[42582] = MEM[35298] + MEM[35377];
assign MEM[42583] = MEM[35299] + MEM[35376];
assign MEM[42584] = MEM[35303] + MEM[35334];
assign MEM[42585] = MEM[35306] + MEM[35374];
assign MEM[42586] = MEM[35308] + MEM[35362];
assign MEM[42587] = MEM[35311] + MEM[35327];
assign MEM[42588] = MEM[35313] + MEM[35373];
assign MEM[42589] = MEM[35314] + MEM[35329];
assign MEM[42590] = MEM[35315] + MEM[35403];
assign MEM[42591] = MEM[35316] + MEM[35333];
assign MEM[42592] = MEM[35318] + MEM[35370];
assign MEM[42593] = MEM[35319] + MEM[35361];
assign MEM[42594] = MEM[35321] + MEM[35328];
assign MEM[42595] = MEM[35324] + MEM[35340];
assign MEM[42596] = MEM[35325] + MEM[35417];
assign MEM[42597] = MEM[35326] + MEM[35379];
assign MEM[42598] = MEM[35331] + MEM[35348];
assign MEM[42599] = MEM[35335] + MEM[35350];
assign MEM[42600] = MEM[35336] + MEM[35398];
assign MEM[42601] = MEM[35337] + MEM[35488];
assign MEM[42602] = MEM[35338] + MEM[35363];
assign MEM[42603] = MEM[35339] + MEM[35394];
assign MEM[42604] = MEM[35341] + MEM[35404];
assign MEM[42605] = MEM[35344] + MEM[35355];
assign MEM[42606] = MEM[35345] + MEM[35445];
assign MEM[42607] = MEM[35351] + MEM[35400];
assign MEM[42608] = MEM[35353] + MEM[35387];
assign MEM[42609] = MEM[35354] + MEM[35424];
assign MEM[42610] = MEM[35360] + MEM[35425];
assign MEM[42611] = MEM[35364] + MEM[35410];
assign MEM[42612] = MEM[35365] + MEM[35455];
assign MEM[42613] = MEM[35366] + MEM[35463];
assign MEM[42614] = MEM[35368] + MEM[35544];
assign MEM[42615] = MEM[35369] + MEM[35401];
assign MEM[42616] = MEM[35371] + MEM[35382];
assign MEM[42617] = MEM[35372] + MEM[35378];
assign MEM[42618] = MEM[35375] + MEM[35477];
assign MEM[42619] = MEM[35380] + MEM[35427];
assign MEM[42620] = MEM[35381] + MEM[35498];
assign MEM[42621] = MEM[35383] + MEM[35441];
assign MEM[42622] = MEM[35384] + MEM[35511];
assign MEM[42623] = MEM[35385] + MEM[35509];
assign MEM[42624] = MEM[35388] + MEM[35413];
assign MEM[42625] = MEM[35389] + MEM[35461];
assign MEM[42626] = MEM[35390] + MEM[35435];
assign MEM[42627] = MEM[35391] + MEM[35490];
assign MEM[42628] = MEM[35392] + MEM[35505];
assign MEM[42629] = MEM[35393] + MEM[35429];
assign MEM[42630] = MEM[35395] + MEM[35432];
assign MEM[42631] = MEM[35397] + MEM[35582];
assign MEM[42632] = MEM[35399] + MEM[35420];
assign MEM[42633] = MEM[35402] + MEM[35520];
assign MEM[42634] = MEM[35405] + MEM[35473];
assign MEM[42635] = MEM[35406] + MEM[35438];
assign MEM[42636] = MEM[35408] + MEM[35568];
assign MEM[42637] = MEM[35409] + MEM[35426];
assign MEM[42638] = MEM[35411] + MEM[35450];
assign MEM[42639] = MEM[35412] + MEM[35479];
assign MEM[42640] = MEM[35414] + MEM[35485];
assign MEM[42641] = MEM[35415] + MEM[35428];
assign MEM[42642] = MEM[35416] + MEM[35439];
assign MEM[42643] = MEM[35418] + MEM[35539];
assign MEM[42644] = MEM[35419] + MEM[35478];
assign MEM[42645] = MEM[35421] + MEM[35458];
assign MEM[42646] = MEM[35422] + MEM[35502];
assign MEM[42647] = MEM[35423] + MEM[35454];
assign MEM[42648] = MEM[35430] + MEM[35487];
assign MEM[42649] = MEM[35431] + MEM[35506];
assign MEM[42650] = MEM[35433] + MEM[35503];
assign MEM[42651] = MEM[35434] + MEM[35468];
assign MEM[42652] = MEM[35436] + MEM[35493];
assign MEM[42653] = MEM[35437] + MEM[35462];
assign MEM[42654] = MEM[35440] + MEM[35459];
assign MEM[42655] = MEM[35442] + MEM[35457];
assign MEM[42656] = MEM[35443] + MEM[35486];
assign MEM[42657] = MEM[35444] + MEM[35500];
assign MEM[42658] = MEM[35446] + MEM[35483];
assign MEM[42659] = MEM[35447] + MEM[35545];
assign MEM[42660] = MEM[35448] + MEM[35489];
assign MEM[42661] = MEM[35449] + MEM[35492];
assign MEM[42662] = MEM[35451] + MEM[35518];
assign MEM[42663] = MEM[35452] + MEM[35541];
assign MEM[42664] = MEM[35456] + MEM[35625];
assign MEM[42665] = MEM[35460] + MEM[35480];
assign MEM[42666] = MEM[35464] + MEM[35475];
assign MEM[42667] = MEM[35465] + MEM[35565];
assign MEM[42668] = MEM[35467] + MEM[35510];
assign MEM[42669] = MEM[35469] + MEM[35525];
assign MEM[42670] = MEM[35470] + MEM[35550];
assign MEM[42671] = MEM[35471] + MEM[35484];
assign MEM[42672] = MEM[35472] + MEM[35549];
assign MEM[42673] = MEM[35474] + MEM[35559];
assign MEM[42674] = MEM[35476] + MEM[35495];
assign MEM[42675] = MEM[35481] + MEM[35583];
assign MEM[42676] = MEM[35482] + MEM[35584];
assign MEM[42677] = MEM[35491] + MEM[35614];
assign MEM[42678] = MEM[35494] + MEM[35530];
assign MEM[42679] = MEM[35496] + MEM[35517];
assign MEM[42680] = MEM[35497] + MEM[35579];
assign MEM[42681] = MEM[35499] + MEM[35571];
assign MEM[42682] = MEM[35501] + MEM[35531];
assign MEM[42683] = MEM[35504] + MEM[35569];
assign MEM[42684] = MEM[35507] + MEM[35566];
assign MEM[42685] = MEM[35508] + MEM[35601];
assign MEM[42686] = MEM[35512] + MEM[35523];
assign MEM[42687] = MEM[35513] + MEM[35540];
assign MEM[42688] = MEM[35514] + MEM[35562];
assign MEM[42689] = MEM[35515] + MEM[35534];
assign MEM[42690] = MEM[35516] + MEM[35546];
assign MEM[42691] = MEM[35519] + MEM[35577];
assign MEM[42692] = MEM[35521] + MEM[35778];
assign MEM[42693] = MEM[35522] + MEM[35661];
assign MEM[42694] = MEM[35524] + MEM[35588];
assign MEM[42695] = MEM[35526] + MEM[35591];
assign MEM[42696] = MEM[35527] + MEM[35597];
assign MEM[42697] = MEM[35528] + MEM[35623];
assign MEM[42698] = MEM[35529] + MEM[35573];
assign MEM[42699] = MEM[35532] + MEM[35557];
assign MEM[42700] = MEM[35533] + MEM[35548];
assign MEM[42701] = MEM[35535] + MEM[35666];
assign MEM[42702] = MEM[35536] + MEM[35592];
assign MEM[42703] = MEM[35537] + MEM[35617];
assign MEM[42704] = MEM[35538] + MEM[35629];
assign MEM[42705] = MEM[35542] + MEM[35632];
assign MEM[42706] = MEM[35543] + MEM[35640];
assign MEM[42707] = MEM[35547] + MEM[35657];
assign MEM[42708] = MEM[35551] + MEM[35558];
assign MEM[42709] = MEM[35552] + MEM[35576];
assign MEM[42710] = MEM[35553] + MEM[35556];
assign MEM[42711] = MEM[35554] + MEM[35590];
assign MEM[42712] = MEM[35555] + MEM[35684];
assign MEM[42713] = MEM[35560] + MEM[35622];
assign MEM[42714] = MEM[35561] + MEM[35641];
assign MEM[42715] = MEM[35563] + MEM[35659];
assign MEM[42716] = MEM[35564] + MEM[35607];
assign MEM[42717] = MEM[35567] + MEM[35616];
assign MEM[42718] = MEM[35570] + MEM[35695];
assign MEM[42719] = MEM[35572] + MEM[35660];
assign MEM[42720] = MEM[35574] + MEM[35693];
assign MEM[42721] = MEM[35575] + MEM[35644];
assign MEM[42722] = MEM[35578] + MEM[35624];
assign MEM[42723] = MEM[35580] + MEM[35630];
assign MEM[42724] = MEM[35581] + MEM[35604];
assign MEM[42725] = MEM[35585] + MEM[35647];
assign MEM[42726] = MEM[35586] + MEM[35593];
assign MEM[42727] = MEM[35587] + MEM[35636];
assign MEM[42728] = MEM[35589] + MEM[35645];
assign MEM[42729] = MEM[35594] + MEM[35687];
assign MEM[42730] = MEM[35595] + MEM[35612];
assign MEM[42731] = MEM[35596] + MEM[35608];
assign MEM[42732] = MEM[35598] + MEM[35733];
assign MEM[42733] = MEM[35599] + MEM[35653];
assign MEM[42734] = MEM[35600] + MEM[35631];
assign MEM[42735] = MEM[35602] + MEM[35682];
assign MEM[42736] = MEM[35603] + MEM[35654];
assign MEM[42737] = MEM[35605] + MEM[35649];
assign MEM[42738] = MEM[35606] + MEM[35658];
assign MEM[42739] = MEM[35609] + MEM[35753];
assign MEM[42740] = MEM[35610] + MEM[35652];
assign MEM[42741] = MEM[35611] + MEM[35795];
assign MEM[42742] = MEM[35613] + MEM[35681];
assign MEM[42743] = MEM[35615] + MEM[35626];
assign MEM[42744] = MEM[35618] + MEM[35664];
assign MEM[42745] = MEM[35619] + MEM[35694];
assign MEM[42746] = MEM[35620] + MEM[35670];
assign MEM[42747] = MEM[35621] + MEM[35705];
assign MEM[42748] = MEM[35627] + MEM[35643];
assign MEM[42749] = MEM[35628] + MEM[35672];
assign MEM[42750] = MEM[35633] + MEM[35714];
assign MEM[42751] = MEM[35634] + MEM[35679];
assign MEM[42752] = MEM[35635] + MEM[35671];
assign MEM[42753] = MEM[35637] + MEM[35692];
assign MEM[42754] = MEM[35638] + MEM[35667];
assign MEM[42755] = MEM[35639] + MEM[35677];
assign MEM[42756] = MEM[35642] + MEM[35669];
assign MEM[42757] = MEM[35646] + MEM[35765];
assign MEM[42758] = MEM[35648] + MEM[35708];
assign MEM[42759] = MEM[35650] + MEM[35697];
assign MEM[42760] = MEM[35651] + MEM[35755];
assign MEM[42761] = MEM[35655] + MEM[35702];
assign MEM[42762] = MEM[35656] + MEM[35691];
assign MEM[42763] = MEM[35662] + MEM[35676];
assign MEM[42764] = MEM[35663] + MEM[35747];
assign MEM[42765] = MEM[35665] + MEM[35875];
assign MEM[42766] = MEM[35668] + MEM[35739];
assign MEM[42767] = MEM[35673] + MEM[35876];
assign MEM[42768] = MEM[35674] + MEM[35763];
assign MEM[42769] = MEM[35675] + MEM[35734];
assign MEM[42770] = MEM[35678] + MEM[35723];
assign MEM[42771] = MEM[35680] + MEM[35743];
assign MEM[42772] = MEM[35683] + MEM[35722];
assign MEM[42773] = MEM[35685] + MEM[35812];
assign MEM[42774] = MEM[35686] + MEM[35793];
assign MEM[42775] = MEM[35688] + MEM[35808];
assign MEM[42776] = MEM[35689] + MEM[35718];
assign MEM[42777] = MEM[35690] + MEM[35696];
assign MEM[42778] = MEM[35698] + MEM[35846];
assign MEM[42779] = MEM[35699] + MEM[35926];
assign MEM[42780] = MEM[35700] + MEM[35716];
assign MEM[42781] = MEM[35701] + MEM[35791];
assign MEM[42782] = MEM[35703] + MEM[35760];
assign MEM[42783] = MEM[35704] + MEM[35726];
assign MEM[42784] = MEM[35706] + MEM[35727];
assign MEM[42785] = MEM[35707] + MEM[35730];
assign MEM[42786] = MEM[35709] + MEM[35786];
assign MEM[42787] = MEM[35710] + MEM[35735];
assign MEM[42788] = MEM[35711] + MEM[35776];
assign MEM[42789] = MEM[35712] + MEM[35737];
assign MEM[42790] = MEM[35713] + MEM[35736];
assign MEM[42791] = MEM[35715] + MEM[35814];
assign MEM[42792] = MEM[35717] + MEM[35877];
assign MEM[42793] = MEM[35719] + MEM[35839];
assign MEM[42794] = MEM[35720] + MEM[35752];
assign MEM[42795] = MEM[35721] + MEM[35804];
assign MEM[42796] = MEM[35724] + MEM[35757];
assign MEM[42797] = MEM[35725] + MEM[35749];
assign MEM[42798] = MEM[35728] + MEM[35887];
assign MEM[42799] = MEM[35729] + MEM[35768];
assign MEM[42800] = MEM[35731] + MEM[35754];
assign MEM[42801] = MEM[35732] + MEM[35785];
assign MEM[42802] = MEM[35738] + MEM[35771];
assign MEM[42803] = MEM[35740] + MEM[35764];
assign MEM[42804] = MEM[35741] + MEM[35794];
assign MEM[42805] = MEM[35742] + MEM[35789];
assign MEM[42806] = MEM[35744] + MEM[35784];
assign MEM[42807] = MEM[35745] + MEM[35820];
assign MEM[42808] = MEM[35746] + MEM[35803];
assign MEM[42809] = MEM[35748] + MEM[35848];
assign MEM[42810] = MEM[35750] + MEM[35833];
assign MEM[42811] = MEM[35751] + MEM[35822];
assign MEM[42812] = MEM[35756] + MEM[35879];
assign MEM[42813] = MEM[35758] + MEM[35866];
assign MEM[42814] = MEM[35759] + MEM[35859];
assign MEM[42815] = MEM[35761] + MEM[35851];
assign MEM[42816] = MEM[35762] + MEM[35817];
assign MEM[42817] = MEM[35766] + MEM[35813];
assign MEM[42818] = MEM[35767] + MEM[35774];
assign MEM[42819] = MEM[35769] + MEM[35816];
assign MEM[42820] = MEM[35770] + MEM[35779];
assign MEM[42821] = MEM[35772] + MEM[35810];
assign MEM[42822] = MEM[35773] + MEM[35811];
assign MEM[42823] = MEM[35775] + MEM[35809];
assign MEM[42824] = MEM[35777] + MEM[35967];
assign MEM[42825] = MEM[35780] + MEM[35838];
assign MEM[42826] = MEM[35781] + MEM[35807];
assign MEM[42827] = MEM[35782] + MEM[35869];
assign MEM[42828] = MEM[35783] + MEM[35871];
assign MEM[42829] = MEM[35787] + MEM[35845];
assign MEM[42830] = MEM[35788] + MEM[35854];
assign MEM[42831] = MEM[35790] + MEM[35819];
assign MEM[42832] = MEM[35792] + MEM[35821];
assign MEM[42833] = MEM[35796] + MEM[35815];
assign MEM[42834] = MEM[35797] + MEM[35832];
assign MEM[42835] = MEM[35798] + MEM[35830];
assign MEM[42836] = MEM[35799] + MEM[36063];
assign MEM[42837] = MEM[35800] + MEM[35825];
assign MEM[42838] = MEM[35801] + MEM[35826];
assign MEM[42839] = MEM[35802] + MEM[35885];
assign MEM[42840] = MEM[35805] + MEM[35849];
assign MEM[42841] = MEM[35806] + MEM[35936];
assign MEM[42842] = MEM[35818] + MEM[35852];
assign MEM[42843] = MEM[35823] + MEM[35893];
assign MEM[42844] = MEM[35824] + MEM[35853];
assign MEM[42845] = MEM[35827] + MEM[35874];
assign MEM[42846] = MEM[35828] + MEM[35873];
assign MEM[42847] = MEM[35829] + MEM[35868];
assign MEM[42848] = MEM[35831] + MEM[35908];
assign MEM[42849] = MEM[35834] + MEM[35939];
assign MEM[42850] = MEM[35835] + MEM[35862];
assign MEM[42851] = MEM[35836] + MEM[35894];
assign MEM[42852] = MEM[35837] + MEM[35855];
assign MEM[42853] = MEM[35840] + MEM[35977];
assign MEM[42854] = MEM[35841] + MEM[35923];
assign MEM[42855] = MEM[35842] + MEM[35941];
assign MEM[42856] = MEM[35843] + MEM[35904];
assign MEM[42857] = MEM[35844] + MEM[35954];
assign MEM[42858] = MEM[35847] + MEM[35872];
assign MEM[42859] = MEM[35850] + MEM[35907];
assign MEM[42860] = MEM[35856] + MEM[35895];
assign MEM[42861] = MEM[35857] + MEM[35930];
assign MEM[42862] = MEM[35858] + MEM[35891];
assign MEM[42863] = MEM[35860] + MEM[35897];
assign MEM[42864] = MEM[35861] + MEM[35963];
assign MEM[42865] = MEM[35863] + MEM[35870];
assign MEM[42866] = MEM[35864] + MEM[35917];
assign MEM[42867] = MEM[35865] + MEM[35937];
assign MEM[42868] = MEM[35867] + MEM[35918];
assign MEM[42869] = MEM[35878] + MEM[36019];
assign MEM[42870] = MEM[35880] + MEM[35900];
assign MEM[42871] = MEM[35881] + MEM[35913];
assign MEM[42872] = MEM[35882] + MEM[35992];
assign MEM[42873] = MEM[35883] + MEM[35911];
assign MEM[42874] = MEM[35884] + MEM[35990];
assign MEM[42875] = MEM[35886] + MEM[35898];
assign MEM[42876] = MEM[35888] + MEM[35905];
assign MEM[42877] = MEM[35889] + MEM[35906];
assign MEM[42878] = MEM[35890] + MEM[35980];
assign MEM[42879] = MEM[35892] + MEM[35986];
assign MEM[42880] = MEM[35896] + MEM[35942];
assign MEM[42881] = MEM[35899] + MEM[35998];
assign MEM[42882] = MEM[35901] + MEM[36043];
assign MEM[42883] = MEM[35902] + MEM[35916];
assign MEM[42884] = MEM[35903] + MEM[36196];
assign MEM[42885] = MEM[35909] + MEM[35966];
assign MEM[42886] = MEM[35910] + MEM[36032];
assign MEM[42887] = MEM[35912] + MEM[35973];
assign MEM[42888] = MEM[35914] + MEM[35948];
assign MEM[42889] = MEM[35915] + MEM[35952];
assign MEM[42890] = MEM[35919] + MEM[36004];
assign MEM[42891] = MEM[35920] + MEM[35991];
assign MEM[42892] = MEM[35921] + MEM[35970];
assign MEM[42893] = MEM[35922] + MEM[35932];
assign MEM[42894] = MEM[35924] + MEM[35983];
assign MEM[42895] = MEM[35925] + MEM[35968];
assign MEM[42896] = MEM[35927] + MEM[35975];
assign MEM[42897] = MEM[35928] + MEM[35951];
assign MEM[42898] = MEM[35929] + MEM[35962];
assign MEM[42899] = MEM[35931] + MEM[35959];
assign MEM[42900] = MEM[35933] + MEM[36084];
assign MEM[42901] = MEM[35934] + MEM[36011];
assign MEM[42902] = MEM[35935] + MEM[35961];
assign MEM[42903] = MEM[35938] + MEM[35969];
assign MEM[42904] = MEM[35940] + MEM[35946];
assign MEM[42905] = MEM[35943] + MEM[36028];
assign MEM[42906] = MEM[35944] + MEM[35999];
assign MEM[42907] = MEM[35945] + MEM[36003];
assign MEM[42908] = MEM[35947] + MEM[35972];
assign MEM[42909] = MEM[35949] + MEM[36020];
assign MEM[42910] = MEM[35950] + MEM[36039];
assign MEM[42911] = MEM[35953] + MEM[36009];
assign MEM[42912] = MEM[35955] + MEM[36005];
assign MEM[42913] = MEM[35956] + MEM[36027];
assign MEM[42914] = MEM[35957] + MEM[36006];
assign MEM[42915] = MEM[35958] + MEM[36010];
assign MEM[42916] = MEM[35960] + MEM[36070];
assign MEM[42917] = MEM[35964] + MEM[36047];
assign MEM[42918] = MEM[35965] + MEM[36051];
assign MEM[42919] = MEM[35971] + MEM[36002];
assign MEM[42920] = MEM[35974] + MEM[36075];
assign MEM[42921] = MEM[35976] + MEM[36012];
assign MEM[42922] = MEM[35978] + MEM[36049];
assign MEM[42923] = MEM[35979] + MEM[36056];
assign MEM[42924] = MEM[35981] + MEM[35987];
assign MEM[42925] = MEM[35982] + MEM[36105];
assign MEM[42926] = MEM[35984] + MEM[36024];
assign MEM[42927] = MEM[35985] + MEM[36031];
assign MEM[42928] = MEM[35988] + MEM[36041];
assign MEM[42929] = MEM[35989] + MEM[36023];
assign MEM[42930] = MEM[35993] + MEM[36030];
assign MEM[42931] = MEM[35994] + MEM[36048];
assign MEM[42932] = MEM[35995] + MEM[36142];
assign MEM[42933] = MEM[35996] + MEM[36037];
assign MEM[42934] = MEM[35997] + MEM[36135];
assign MEM[42935] = MEM[36000] + MEM[36038];
assign MEM[42936] = MEM[36001] + MEM[36061];
assign MEM[42937] = MEM[36007] + MEM[36046];
assign MEM[42938] = MEM[36008] + MEM[36050];
assign MEM[42939] = MEM[36013] + MEM[36121];
assign MEM[42940] = MEM[36014] + MEM[36055];
assign MEM[42941] = MEM[36015] + MEM[36108];
assign MEM[42942] = MEM[36016] + MEM[36111];
assign MEM[42943] = MEM[36017] + MEM[36036];
assign MEM[42944] = MEM[36018] + MEM[36058];
assign MEM[42945] = MEM[36021] + MEM[36217];
assign MEM[42946] = MEM[36022] + MEM[36148];
assign MEM[42947] = MEM[36025] + MEM[36190];
assign MEM[42948] = MEM[36026] + MEM[36091];
assign MEM[42949] = MEM[36029] + MEM[36062];
assign MEM[42950] = MEM[36033] + MEM[36141];
assign MEM[42951] = MEM[36034] + MEM[36080];
assign MEM[42952] = MEM[36035] + MEM[36103];
assign MEM[42953] = MEM[36040] + MEM[36116];
assign MEM[42954] = MEM[36042] + MEM[36101];
assign MEM[42955] = MEM[36044] + MEM[36092];
assign MEM[42956] = MEM[36045] + MEM[36064];
assign MEM[42957] = MEM[36052] + MEM[36066];
assign MEM[42958] = MEM[36053] + MEM[36089];
assign MEM[42959] = MEM[36054] + MEM[36107];
assign MEM[42960] = MEM[36057] + MEM[36069];
assign MEM[42961] = MEM[36059] + MEM[36128];
assign MEM[42962] = MEM[36060] + MEM[36109];
assign MEM[42963] = MEM[36065] + MEM[36255];
assign MEM[42964] = MEM[36067] + MEM[36072];
assign MEM[42965] = MEM[36068] + MEM[36078];
assign MEM[42966] = MEM[36071] + MEM[36131];
assign MEM[42967] = MEM[36073] + MEM[36117];
assign MEM[42968] = MEM[36074] + MEM[36178];
assign MEM[42969] = MEM[36076] + MEM[36153];
assign MEM[42970] = MEM[36077] + MEM[36173];
assign MEM[42971] = MEM[36079] + MEM[36209];
assign MEM[42972] = MEM[36081] + MEM[36134];
assign MEM[42973] = MEM[36082] + MEM[36225];
assign MEM[42974] = MEM[36083] + MEM[36106];
assign MEM[42975] = MEM[36085] + MEM[36157];
assign MEM[42976] = MEM[36086] + MEM[36100];
assign MEM[42977] = MEM[36087] + MEM[36177];
assign MEM[42978] = MEM[36088] + MEM[36114];
assign MEM[42979] = MEM[36090] + MEM[36214];
assign MEM[42980] = MEM[36093] + MEM[36175];
assign MEM[42981] = MEM[36094] + MEM[36144];
assign MEM[42982] = MEM[36095] + MEM[36137];
assign MEM[42983] = MEM[36096] + MEM[36158];
assign MEM[42984] = MEM[36097] + MEM[36136];
assign MEM[42985] = MEM[36098] + MEM[36110];
assign MEM[42986] = MEM[36099] + MEM[36124];
assign MEM[42987] = MEM[36102] + MEM[36268];
assign MEM[42988] = MEM[36104] + MEM[36119];
assign MEM[42989] = MEM[36112] + MEM[36169];
assign MEM[42990] = MEM[36113] + MEM[36149];
assign MEM[42991] = MEM[36115] + MEM[36143];
assign MEM[42992] = MEM[36118] + MEM[36170];
assign MEM[42993] = MEM[36120] + MEM[36219];
assign MEM[42994] = MEM[36122] + MEM[36204];
assign MEM[42995] = MEM[36123] + MEM[36226];
assign MEM[42996] = MEM[36125] + MEM[36192];
assign MEM[42997] = MEM[36126] + MEM[36185];
assign MEM[42998] = MEM[36127] + MEM[36172];
assign MEM[42999] = MEM[36129] + MEM[36156];
assign MEM[43000] = MEM[36130] + MEM[36212];
assign MEM[43001] = MEM[36132] + MEM[36145];
assign MEM[43002] = MEM[36133] + MEM[36171];
assign MEM[43003] = MEM[36138] + MEM[36248];
assign MEM[43004] = MEM[36139] + MEM[36200];
assign MEM[43005] = MEM[36140] + MEM[36315];
assign MEM[43006] = MEM[36146] + MEM[36161];
assign MEM[43007] = MEM[36147] + MEM[36180];
assign MEM[43008] = MEM[36150] + MEM[36174];
assign MEM[43009] = MEM[36151] + MEM[36198];
assign MEM[43010] = MEM[36152] + MEM[36179];
assign MEM[43011] = MEM[36154] + MEM[36202];
assign MEM[43012] = MEM[36155] + MEM[36238];
assign MEM[43013] = MEM[36159] + MEM[36272];
assign MEM[43014] = MEM[36160] + MEM[36197];
assign MEM[43015] = MEM[36162] + MEM[36241];
assign MEM[43016] = MEM[36163] + MEM[36257];
assign MEM[43017] = MEM[36164] + MEM[36176];
assign MEM[43018] = MEM[36165] + MEM[36222];
assign MEM[43019] = MEM[36166] + MEM[36201];
assign MEM[43020] = MEM[36167] + MEM[36262];
assign MEM[43021] = MEM[36168] + MEM[36213];
assign MEM[43022] = MEM[36181] + MEM[36321];
assign MEM[43023] = MEM[36182] + MEM[36211];
assign MEM[43024] = MEM[36183] + MEM[36249];
assign MEM[43025] = MEM[36184] + MEM[36231];
assign MEM[43026] = MEM[36186] + MEM[36210];
assign MEM[43027] = MEM[36187] + MEM[36220];
assign MEM[43028] = MEM[36188] + MEM[36264];
assign MEM[43029] = MEM[36189] + MEM[36215];
assign MEM[43030] = MEM[36191] + MEM[36273];
assign MEM[43031] = MEM[36193] + MEM[36260];
assign MEM[43032] = MEM[36194] + MEM[36252];
assign MEM[43033] = MEM[36195] + MEM[36288];
assign MEM[43034] = MEM[36199] + MEM[36240];
assign MEM[43035] = MEM[36203] + MEM[36459];
assign MEM[43036] = MEM[36205] + MEM[36256];
assign MEM[43037] = MEM[36206] + MEM[36293];
assign MEM[43038] = MEM[36207] + MEM[36305];
assign MEM[43039] = MEM[36208] + MEM[36228];
assign MEM[43040] = MEM[36216] + MEM[36300];
assign MEM[43041] = MEM[36218] + MEM[36266];
assign MEM[43042] = MEM[36221] + MEM[36276];
assign MEM[43043] = MEM[36223] + MEM[36244];
assign MEM[43044] = MEM[36224] + MEM[36233];
assign MEM[43045] = MEM[36227] + MEM[36325];
assign MEM[43046] = MEM[36229] + MEM[36360];
assign MEM[43047] = MEM[36230] + MEM[36261];
assign MEM[43048] = MEM[36232] + MEM[36322];
assign MEM[43049] = MEM[36234] + MEM[36250];
assign MEM[43050] = MEM[36235] + MEM[36287];
assign MEM[43051] = MEM[36236] + MEM[36277];
assign MEM[43052] = MEM[36237] + MEM[36259];
assign MEM[43053] = MEM[36239] + MEM[36283];
assign MEM[43054] = MEM[36242] + MEM[36312];
assign MEM[43055] = MEM[36243] + MEM[36331];
assign MEM[43056] = MEM[36245] + MEM[36278];
assign MEM[43057] = MEM[36246] + MEM[36341];
assign MEM[43058] = MEM[36247] + MEM[36289];
assign MEM[43059] = MEM[36251] + MEM[36274];
assign MEM[43060] = MEM[36253] + MEM[36269];
assign MEM[43061] = MEM[36254] + MEM[36281];
assign MEM[43062] = MEM[36258] + MEM[36329];
assign MEM[43063] = MEM[36263] + MEM[36396];
assign MEM[43064] = MEM[36265] + MEM[36299];
assign MEM[43065] = MEM[36267] + MEM[36357];
assign MEM[43066] = MEM[36270] + MEM[36422];
assign MEM[43067] = MEM[36271] + MEM[36372];
assign MEM[43068] = MEM[36275] + MEM[36318];
assign MEM[43069] = MEM[36279] + MEM[36367];
assign MEM[43070] = MEM[36280] + MEM[36292];
assign MEM[43071] = MEM[36282] + MEM[36333];
assign MEM[43072] = MEM[36284] + MEM[36296];
assign MEM[43073] = MEM[36285] + MEM[36416];
assign MEM[43074] = MEM[36286] + MEM[36429];
assign MEM[43075] = MEM[36290] + MEM[36356];
assign MEM[43076] = MEM[36291] + MEM[36380];
assign MEM[43077] = MEM[36294] + MEM[36307];
assign MEM[43078] = MEM[36295] + MEM[36382];
assign MEM[43079] = MEM[36297] + MEM[36427];
assign MEM[43080] = MEM[36298] + MEM[36399];
assign MEM[43081] = MEM[36301] + MEM[36347];
assign MEM[43082] = MEM[36302] + MEM[36345];
assign MEM[43083] = MEM[36303] + MEM[36311];
assign MEM[43084] = MEM[36304] + MEM[36391];
assign MEM[43085] = MEM[36306] + MEM[36335];
assign MEM[43086] = MEM[36308] + MEM[36395];
assign MEM[43087] = MEM[36309] + MEM[36420];
assign MEM[43088] = MEM[36310] + MEM[36417];
assign MEM[43089] = MEM[36313] + MEM[36343];
assign MEM[43090] = MEM[36314] + MEM[36415];
assign MEM[43091] = MEM[36316] + MEM[36330];
assign MEM[43092] = MEM[36317] + MEM[36531];
assign MEM[43093] = MEM[36319] + MEM[36358];
assign MEM[43094] = MEM[36320] + MEM[36406];
assign MEM[43095] = MEM[36323] + MEM[36379];
assign MEM[43096] = MEM[36324] + MEM[36328];
assign MEM[43097] = MEM[36326] + MEM[36410];
assign MEM[43098] = MEM[36327] + MEM[36378];
assign MEM[43099] = MEM[36332] + MEM[36403];
assign MEM[43100] = MEM[36334] + MEM[36404];
assign MEM[43101] = MEM[36336] + MEM[36377];
assign MEM[43102] = MEM[36337] + MEM[36411];
assign MEM[43103] = MEM[36338] + MEM[36408];
assign MEM[43104] = MEM[36339] + MEM[36374];
assign MEM[43105] = MEM[36340] + MEM[36381];
assign MEM[43106] = MEM[36342] + MEM[36419];
assign MEM[43107] = MEM[36344] + MEM[36373];
assign MEM[43108] = MEM[36346] + MEM[36363];
assign MEM[43109] = MEM[36348] + MEM[36393];
assign MEM[43110] = MEM[36349] + MEM[36375];
assign MEM[43111] = MEM[36350] + MEM[36366];
assign MEM[43112] = MEM[36351] + MEM[36392];
assign MEM[43113] = MEM[36352] + MEM[36431];
assign MEM[43114] = MEM[36353] + MEM[36370];
assign MEM[43115] = MEM[36354] + MEM[36394];
assign MEM[43116] = MEM[36355] + MEM[36440];
assign MEM[43117] = MEM[36359] + MEM[36390];
assign MEM[43118] = MEM[36361] + MEM[36405];
assign MEM[43119] = MEM[36362] + MEM[36452];
assign MEM[43120] = MEM[36364] + MEM[36389];
assign MEM[43121] = MEM[36365] + MEM[36397];
assign MEM[43122] = MEM[36368] + MEM[36402];
assign MEM[43123] = MEM[36369] + MEM[36438];
assign MEM[43124] = MEM[36371] + MEM[36407];
assign MEM[43125] = MEM[36376] + MEM[36435];
assign MEM[43126] = MEM[36383] + MEM[36451];
assign MEM[43127] = MEM[36384] + MEM[36439];
assign MEM[43128] = MEM[36385] + MEM[36475];
assign MEM[43129] = MEM[36386] + MEM[36460];
assign MEM[43130] = MEM[36387] + MEM[36483];
assign MEM[43131] = MEM[36388] + MEM[36423];
assign MEM[43132] = MEM[36398] + MEM[36432];
assign MEM[43133] = MEM[36400] + MEM[36447];
assign MEM[43134] = MEM[36401] + MEM[36433];
assign MEM[43135] = MEM[36409] + MEM[36584];
assign MEM[43136] = MEM[36412] + MEM[36546];
assign MEM[43137] = MEM[36413] + MEM[36477];
assign MEM[43138] = MEM[36414] + MEM[36480];
assign MEM[43139] = MEM[36418] + MEM[36466];
assign MEM[43140] = MEM[36421] + MEM[36576];
assign MEM[43141] = MEM[36424] + MEM[36484];
assign MEM[43142] = MEM[36425] + MEM[36497];
assign MEM[43143] = MEM[36426] + MEM[36479];
assign MEM[43144] = MEM[36428] + MEM[36478];
assign MEM[43145] = MEM[36430] + MEM[36472];
assign MEM[43146] = MEM[36434] + MEM[36555];
assign MEM[43147] = MEM[36436] + MEM[36572];
assign MEM[43148] = MEM[36437] + MEM[36445];
assign MEM[43149] = MEM[36441] + MEM[36474];
assign MEM[43150] = MEM[36442] + MEM[36505];
assign MEM[43151] = MEM[36443] + MEM[36490];
assign MEM[43152] = MEM[36444] + MEM[36487];
assign MEM[43153] = MEM[36446] + MEM[36455];
assign MEM[43154] = MEM[36448] + MEM[36463];
assign MEM[43155] = MEM[36449] + MEM[36575];
assign MEM[43156] = MEM[36450] + MEM[36522];
assign MEM[43157] = MEM[36453] + MEM[36500];
assign MEM[43158] = MEM[36454] + MEM[36504];
assign MEM[43159] = MEM[36456] + MEM[36697];
assign MEM[43160] = MEM[36457] + MEM[36561];
assign MEM[43161] = MEM[36458] + MEM[36517];
assign MEM[43162] = MEM[36461] + MEM[36467];
assign MEM[43163] = MEM[36462] + MEM[36527];
assign MEM[43164] = MEM[36464] + MEM[36537];
assign MEM[43165] = MEM[36465] + MEM[36548];
assign MEM[43166] = MEM[36468] + MEM[36544];
assign MEM[43167] = MEM[36469] + MEM[36526];
assign MEM[43168] = MEM[36470] + MEM[36509];
assign MEM[43169] = MEM[36471] + MEM[36503];
assign MEM[43170] = MEM[36473] + MEM[36562];
assign MEM[43171] = MEM[36476] + MEM[36543];
assign MEM[43172] = MEM[36481] + MEM[36494];
assign MEM[43173] = MEM[36482] + MEM[36559];
assign MEM[43174] = MEM[36485] + MEM[36563];
assign MEM[43175] = MEM[36486] + MEM[36523];
assign MEM[43176] = MEM[36488] + MEM[36520];
assign MEM[43177] = MEM[36489] + MEM[36627];
assign MEM[43178] = MEM[36491] + MEM[36525];
assign MEM[43179] = MEM[36492] + MEM[36499];
assign MEM[43180] = MEM[36493] + MEM[36621];
assign MEM[43181] = MEM[36495] + MEM[36579];
assign MEM[43182] = MEM[36496] + MEM[36626];
assign MEM[43183] = MEM[36498] + MEM[36506];
assign MEM[43184] = MEM[36501] + MEM[36588];
assign MEM[43185] = MEM[36502] + MEM[36512];
assign MEM[43186] = MEM[36507] + MEM[36552];
assign MEM[43187] = MEM[36508] + MEM[36536];
assign MEM[43188] = MEM[36510] + MEM[36597];
assign MEM[43189] = MEM[36511] + MEM[36640];
assign MEM[43190] = MEM[36513] + MEM[36530];
assign MEM[43191] = MEM[36514] + MEM[36587];
assign MEM[43192] = MEM[36515] + MEM[36592];
assign MEM[43193] = MEM[36516] + MEM[36569];
assign MEM[43194] = MEM[36518] + MEM[36655];
assign MEM[43195] = MEM[36519] + MEM[36591];
assign MEM[43196] = MEM[36521] + MEM[36553];
assign MEM[43197] = MEM[36524] + MEM[36702];
assign MEM[43198] = MEM[36528] + MEM[36586];
assign MEM[43199] = MEM[36529] + MEM[36534];
assign MEM[43200] = MEM[36532] + MEM[36565];
assign MEM[43201] = MEM[36533] + MEM[36620];
assign MEM[43202] = MEM[36535] + MEM[36570];
assign MEM[43203] = MEM[36538] + MEM[36577];
assign MEM[43204] = MEM[36539] + MEM[36571];
assign MEM[43205] = MEM[36540] + MEM[36568];
assign MEM[43206] = MEM[36541] + MEM[36551];
assign MEM[43207] = MEM[36542] + MEM[36638];
assign MEM[43208] = MEM[36545] + MEM[36645];
assign MEM[43209] = MEM[36547] + MEM[36573];
assign MEM[43210] = MEM[36549] + MEM[36560];
assign MEM[43211] = MEM[36550] + MEM[36578];
assign MEM[43212] = MEM[36554] + MEM[36582];
assign MEM[43213] = MEM[36556] + MEM[36631];
assign MEM[43214] = MEM[36557] + MEM[36658];
assign MEM[43215] = MEM[36558] + MEM[36585];
assign MEM[43216] = MEM[36564] + MEM[36601];
assign MEM[43217] = MEM[36566] + MEM[36704];
assign MEM[43218] = MEM[36567] + MEM[36624];
assign MEM[43219] = MEM[36574] + MEM[36644];
assign MEM[43220] = MEM[36580] + MEM[36623];
assign MEM[43221] = MEM[36581] + MEM[36602];
assign MEM[43222] = MEM[36583] + MEM[36636];
assign MEM[43223] = MEM[36589] + MEM[36670];
assign MEM[43224] = MEM[36590] + MEM[36666];
assign MEM[43225] = MEM[36593] + MEM[36660];
assign MEM[43226] = MEM[36594] + MEM[36651];
assign MEM[43227] = MEM[36595] + MEM[36647];
assign MEM[43228] = MEM[36596] + MEM[36824];
assign MEM[43229] = MEM[36598] + MEM[36608];
assign MEM[43230] = MEM[36599] + MEM[36612];
assign MEM[43231] = MEM[36600] + MEM[36606];
assign MEM[43232] = MEM[36603] + MEM[36667];
assign MEM[43233] = MEM[36604] + MEM[36690];
assign MEM[43234] = MEM[36605] + MEM[36628];
assign MEM[43235] = MEM[36607] + MEM[36805];
assign MEM[43236] = MEM[36609] + MEM[36686];
assign MEM[43237] = MEM[36610] + MEM[36694];
assign MEM[43238] = MEM[36611] + MEM[36688];
assign MEM[43239] = MEM[36613] + MEM[36659];
assign MEM[43240] = MEM[36614] + MEM[36632];
assign MEM[43241] = MEM[36615] + MEM[36662];
assign MEM[43242] = MEM[36616] + MEM[36689];
assign MEM[43243] = MEM[36617] + MEM[36641];
assign MEM[43244] = MEM[36618] + MEM[36733];
assign MEM[43245] = MEM[36619] + MEM[36652];
assign MEM[43246] = MEM[36622] + MEM[36687];
assign MEM[43247] = MEM[36625] + MEM[36635];
assign MEM[43248] = MEM[36629] + MEM[36823];
assign MEM[43249] = MEM[36630] + MEM[36634];
assign MEM[43250] = MEM[36633] + MEM[36654];
assign MEM[43251] = MEM[36637] + MEM[36755];
assign MEM[43252] = MEM[36639] + MEM[36668];
assign MEM[43253] = MEM[36642] + MEM[36677];
assign MEM[43254] = MEM[36643] + MEM[36676];
assign MEM[43255] = MEM[36646] + MEM[36737];
assign MEM[43256] = MEM[36648] + MEM[36729];
assign MEM[43257] = MEM[36649] + MEM[36650];
assign MEM[43258] = MEM[36653] + MEM[36709];
assign MEM[43259] = MEM[36656] + MEM[36724];
assign MEM[43260] = MEM[36657] + MEM[36713];
assign MEM[43261] = MEM[36661] + MEM[36749];
assign MEM[43262] = MEM[36663] + MEM[36740];
assign MEM[43263] = MEM[36664] + MEM[36760];
assign MEM[43264] = MEM[36665] + MEM[36714];
assign MEM[43265] = MEM[36669] + MEM[36691];
assign MEM[43266] = MEM[36671] + MEM[36678];
assign MEM[43267] = MEM[36672] + MEM[36710];
assign MEM[43268] = MEM[36673] + MEM[36807];
assign MEM[43269] = MEM[36674] + MEM[36763];
assign MEM[43270] = MEM[36675] + MEM[36700];
assign MEM[43271] = MEM[36679] + MEM[36793];
assign MEM[43272] = MEM[36680] + MEM[36703];
assign MEM[43273] = MEM[36681] + MEM[36730];
assign MEM[43274] = MEM[36682] + MEM[36695];
assign MEM[43275] = MEM[36683] + MEM[36701];
assign MEM[43276] = MEM[36684] + MEM[36762];
assign MEM[43277] = MEM[36685] + MEM[36829];
assign MEM[43278] = MEM[36692] + MEM[36725];
assign MEM[43279] = MEM[36693] + MEM[36708];
assign MEM[43280] = MEM[36696] + MEM[36735];
assign MEM[43281] = MEM[36698] + MEM[36723];
assign MEM[43282] = MEM[36699] + MEM[36817];
assign MEM[43283] = MEM[36705] + MEM[36711];
assign MEM[43284] = MEM[36706] + MEM[36743];
assign MEM[43285] = MEM[36707] + MEM[36719];
assign MEM[43286] = MEM[36712] + MEM[36739];
assign MEM[43287] = MEM[36715] + MEM[36776];
assign MEM[43288] = MEM[36716] + MEM[36750];
assign MEM[43289] = MEM[36717] + MEM[36771];
assign MEM[43290] = MEM[36718] + MEM[36780];
assign MEM[43291] = MEM[36720] + MEM[36752];
assign MEM[43292] = MEM[36721] + MEM[36732];
assign MEM[43293] = MEM[36722] + MEM[36827];
assign MEM[43294] = MEM[36726] + MEM[36789];
assign MEM[43295] = MEM[36727] + MEM[36779];
assign MEM[43296] = MEM[36728] + MEM[36754];
assign MEM[43297] = MEM[36731] + MEM[36803];
assign MEM[43298] = MEM[36734] + MEM[36873];
assign MEM[43299] = MEM[36736] + MEM[36865];
assign MEM[43300] = MEM[36738] + MEM[36769];
assign MEM[43301] = MEM[36741] + MEM[36778];
assign MEM[43302] = MEM[36742] + MEM[36809];
assign MEM[43303] = MEM[36744] + MEM[36821];
assign MEM[43304] = MEM[36745] + MEM[36781];
assign MEM[43305] = MEM[36746] + MEM[36772];
assign MEM[43306] = MEM[36747] + MEM[36839];
assign MEM[43307] = MEM[36748] + MEM[36757];
assign MEM[43308] = MEM[36751] + MEM[36777];
assign MEM[43309] = MEM[36753] + MEM[36795];
assign MEM[43310] = MEM[36756] + MEM[36888];
assign MEM[43311] = MEM[36758] + MEM[36878];
assign MEM[43312] = MEM[36759] + MEM[36775];
assign MEM[43313] = MEM[36761] + MEM[36810];
assign MEM[43314] = MEM[36764] + MEM[36846];
assign MEM[43315] = MEM[36765] + MEM[36826];
assign MEM[43316] = MEM[36766] + MEM[36782];
assign MEM[43317] = MEM[36767] + MEM[36863];
assign MEM[43318] = MEM[36768] + MEM[36843];
assign MEM[43319] = MEM[36770] + MEM[36783];
assign MEM[43320] = MEM[36773] + MEM[36830];
assign MEM[43321] = MEM[36774] + MEM[36798];
assign MEM[43322] = MEM[36784] + MEM[36901];
assign MEM[43323] = MEM[36785] + MEM[36853];
assign MEM[43324] = MEM[36786] + MEM[36818];
assign MEM[43325] = MEM[36787] + MEM[36910];
assign MEM[43326] = MEM[36788] + MEM[36811];
assign MEM[43327] = MEM[36790] + MEM[36849];
assign MEM[43328] = MEM[36791] + MEM[36801];
assign MEM[43329] = MEM[36792] + MEM[36820];
assign MEM[43330] = MEM[36794] + MEM[36914];
assign MEM[43331] = MEM[36796] + MEM[36831];
assign MEM[43332] = MEM[36797] + MEM[36834];
assign MEM[43333] = MEM[36799] + MEM[36847];
assign MEM[43334] = MEM[36800] + MEM[36837];
assign MEM[43335] = MEM[36802] + MEM[36893];
assign MEM[43336] = MEM[36804] + MEM[36838];
assign MEM[43337] = MEM[36806] + MEM[36933];
assign MEM[43338] = MEM[36808] + MEM[36859];
assign MEM[43339] = MEM[36812] + MEM[36879];
assign MEM[43340] = MEM[36813] + MEM[36898];
assign MEM[43341] = MEM[36814] + MEM[36972];
assign MEM[43342] = MEM[36815] + MEM[36897];
assign MEM[43343] = MEM[36816] + MEM[36877];
assign MEM[43344] = MEM[36819] + MEM[36855];
assign MEM[43345] = MEM[36822] + MEM[36866];
assign MEM[43346] = MEM[36825] + MEM[36884];
assign MEM[43347] = MEM[36828] + MEM[36976];
assign MEM[43348] = MEM[36832] + MEM[36858];
assign MEM[43349] = MEM[36833] + MEM[36852];
assign MEM[43350] = MEM[36835] + MEM[36890];
assign MEM[43351] = MEM[36836] + MEM[36875];
assign MEM[43352] = MEM[36840] + MEM[36864];
assign MEM[43353] = MEM[36841] + MEM[36899];
assign MEM[43354] = MEM[36842] + MEM[36924];
assign MEM[43355] = MEM[36844] + MEM[36915];
assign MEM[43356] = MEM[36845] + MEM[36848];
assign MEM[43357] = MEM[36850] + MEM[36880];
assign MEM[43358] = MEM[36851] + MEM[36896];
assign MEM[43359] = MEM[36854] + MEM[36870];
assign MEM[43360] = MEM[36856] + MEM[36894];
assign MEM[43361] = MEM[36857] + MEM[36928];
assign MEM[43362] = MEM[36860] + MEM[36961];
assign MEM[43363] = MEM[36861] + MEM[36934];
assign MEM[43364] = MEM[36862] + MEM[36867];
assign MEM[43365] = MEM[36868] + MEM[36886];
assign MEM[43366] = MEM[36869] + MEM[36968];
assign MEM[43367] = MEM[36871] + MEM[36882];
assign MEM[43368] = MEM[36872] + MEM[36935];
assign MEM[43369] = MEM[36874] + MEM[36959];
assign MEM[43370] = MEM[36876] + MEM[36908];
assign MEM[43371] = MEM[36881] + MEM[36975];
assign MEM[43372] = MEM[36883] + MEM[36909];
assign MEM[43373] = MEM[36885] + MEM[36907];
assign MEM[43374] = MEM[36887] + MEM[36923];
assign MEM[43375] = MEM[36889] + MEM[36917];
assign MEM[43376] = MEM[36891] + MEM[37032];
assign MEM[43377] = MEM[36892] + MEM[36939];
assign MEM[43378] = MEM[36895] + MEM[36922];
assign MEM[43379] = MEM[36900] + MEM[36950];
assign MEM[43380] = MEM[36902] + MEM[36920];
assign MEM[43381] = MEM[36903] + MEM[36988];
assign MEM[43382] = MEM[36904] + MEM[36919];
assign MEM[43383] = MEM[36905] + MEM[36918];
assign MEM[43384] = MEM[36906] + MEM[36940];
assign MEM[43385] = MEM[36911] + MEM[36982];
assign MEM[43386] = MEM[36912] + MEM[37075];
assign MEM[43387] = MEM[36913] + MEM[37010];
assign MEM[43388] = MEM[36916] + MEM[36962];
assign MEM[43389] = MEM[36921] + MEM[36960];
assign MEM[43390] = MEM[36925] + MEM[37008];
assign MEM[43391] = MEM[36926] + MEM[37053];
assign MEM[43392] = MEM[36927] + MEM[36977];
assign MEM[43393] = MEM[36929] + MEM[36952];
assign MEM[43394] = MEM[36930] + MEM[36948];
assign MEM[43395] = MEM[36931] + MEM[36991];
assign MEM[43396] = MEM[36932] + MEM[37031];
assign MEM[43397] = MEM[36936] + MEM[36994];
assign MEM[43398] = MEM[36937] + MEM[36979];
assign MEM[43399] = MEM[36938] + MEM[36985];
assign MEM[43400] = MEM[36941] + MEM[36998];
assign MEM[43401] = MEM[36942] + MEM[36970];
assign MEM[43402] = MEM[36943] + MEM[36944];
assign MEM[43403] = MEM[36945] + MEM[37040];
assign MEM[43404] = MEM[36946] + MEM[36971];
assign MEM[43405] = MEM[36947] + MEM[37024];
assign MEM[43406] = MEM[36949] + MEM[37005];
assign MEM[43407] = MEM[36951] + MEM[36966];
assign MEM[43408] = MEM[36953] + MEM[36958];
assign MEM[43409] = MEM[36954] + MEM[37023];
assign MEM[43410] = MEM[36955] + MEM[37079];
assign MEM[43411] = MEM[36956] + MEM[37014];
assign MEM[43412] = MEM[36957] + MEM[37052];
assign MEM[43413] = MEM[36963] + MEM[37020];
assign MEM[43414] = MEM[36964] + MEM[36986];
assign MEM[43415] = MEM[36965] + MEM[37041];
assign MEM[43416] = MEM[36967] + MEM[37126];
assign MEM[43417] = MEM[36969] + MEM[37007];
assign MEM[43418] = MEM[36973] + MEM[37006];
assign MEM[43419] = MEM[36974] + MEM[37057];
assign MEM[43420] = MEM[36978] + MEM[37013];
assign MEM[43421] = MEM[36980] + MEM[37018];
assign MEM[43422] = MEM[36981] + MEM[37004];
assign MEM[43423] = MEM[36983] + MEM[37162];
assign MEM[43424] = MEM[36984] + MEM[37066];
assign MEM[43425] = MEM[36987] + MEM[37071];
assign MEM[43426] = MEM[36989] + MEM[37026];
assign MEM[43427] = MEM[36990] + MEM[37034];
assign MEM[43428] = MEM[36992] + MEM[37171];
assign MEM[43429] = MEM[36993] + MEM[36997];
assign MEM[43430] = MEM[36995] + MEM[37077];
assign MEM[43431] = MEM[36996] + MEM[37042];
assign MEM[43432] = MEM[36999] + MEM[37086];
assign MEM[43433] = MEM[37000] + MEM[37029];
assign MEM[43434] = MEM[37001] + MEM[37129];
assign MEM[43435] = MEM[37002] + MEM[37098];
assign MEM[43436] = MEM[37003] + MEM[37060];
assign MEM[43437] = MEM[37009] + MEM[37045];
assign MEM[43438] = MEM[37011] + MEM[37028];
assign MEM[43439] = MEM[37012] + MEM[37058];
assign MEM[43440] = MEM[37015] + MEM[37049];
assign MEM[43441] = MEM[37016] + MEM[37050];
assign MEM[43442] = MEM[37017] + MEM[37124];
assign MEM[43443] = MEM[37019] + MEM[37165];
assign MEM[43444] = MEM[37021] + MEM[37096];
assign MEM[43445] = MEM[37022] + MEM[37046];
assign MEM[43446] = MEM[37025] + MEM[37103];
assign MEM[43447] = MEM[37027] + MEM[37087];
assign MEM[43448] = MEM[37030] + MEM[37189];
assign MEM[43449] = MEM[37033] + MEM[37173];
assign MEM[43450] = MEM[37035] + MEM[37155];
assign MEM[43451] = MEM[37036] + MEM[37151];
assign MEM[43452] = MEM[37037] + MEM[37056];
assign MEM[43453] = MEM[37038] + MEM[37188];
assign MEM[43454] = MEM[37039] + MEM[37084];
assign MEM[43455] = MEM[37043] + MEM[37068];
assign MEM[43456] = MEM[37044] + MEM[37117];
assign MEM[43457] = MEM[37047] + MEM[37061];
assign MEM[43458] = MEM[37048] + MEM[37102];
assign MEM[43459] = MEM[37051] + MEM[37081];
assign MEM[43460] = MEM[37054] + MEM[37065];
assign MEM[43461] = MEM[37055] + MEM[37125];
assign MEM[43462] = MEM[37059] + MEM[37069];
assign MEM[43463] = MEM[37062] + MEM[37115];
assign MEM[43464] = MEM[37063] + MEM[37148];
assign MEM[43465] = MEM[37064] + MEM[37223];
assign MEM[43466] = MEM[37067] + MEM[37109];
assign MEM[43467] = MEM[37070] + MEM[37242];
assign MEM[43468] = MEM[37072] + MEM[37090];
assign MEM[43469] = MEM[37073] + MEM[37132];
assign MEM[43470] = MEM[37074] + MEM[37135];
assign MEM[43471] = MEM[37076] + MEM[37232];
assign MEM[43472] = MEM[37078] + MEM[37105];
assign MEM[43473] = MEM[37080] + MEM[37123];
assign MEM[43474] = MEM[37082] + MEM[37094];
assign MEM[43475] = MEM[37083] + MEM[37101];
assign MEM[43476] = MEM[37085] + MEM[37133];
assign MEM[43477] = MEM[37088] + MEM[37119];
assign MEM[43478] = MEM[37089] + MEM[37131];
assign MEM[43479] = MEM[37091] + MEM[37140];
assign MEM[43480] = MEM[37092] + MEM[37099];
assign MEM[43481] = MEM[37093] + MEM[37100];
assign MEM[43482] = MEM[37095] + MEM[37246];
assign MEM[43483] = MEM[37097] + MEM[37179];
assign MEM[43484] = MEM[37104] + MEM[37138];
assign MEM[43485] = MEM[37106] + MEM[37145];
assign MEM[43486] = MEM[37107] + MEM[37214];
assign MEM[43487] = MEM[37108] + MEM[37118];
assign MEM[43488] = MEM[37110] + MEM[37120];
assign MEM[43489] = MEM[37111] + MEM[37227];
assign MEM[43490] = MEM[37112] + MEM[37128];
assign MEM[43491] = MEM[37113] + MEM[37238];
assign MEM[43492] = MEM[37114] + MEM[37326];
assign MEM[43493] = MEM[37116] + MEM[37184];
assign MEM[43494] = MEM[37121] + MEM[37136];
assign MEM[43495] = MEM[37122] + MEM[37159];
assign MEM[43496] = MEM[37127] + MEM[37150];
assign MEM[43497] = MEM[37130] + MEM[37289];
assign MEM[43498] = MEM[37134] + MEM[37257];
assign MEM[43499] = MEM[37137] + MEM[37201];
assign MEM[43500] = MEM[37139] + MEM[37191];
assign MEM[43501] = MEM[37141] + MEM[37241];
assign MEM[43502] = MEM[37142] + MEM[37198];
assign MEM[43503] = MEM[37143] + MEM[37182];
assign MEM[43504] = MEM[37144] + MEM[37157];
assign MEM[43505] = MEM[37146] + MEM[37211];
assign MEM[43506] = MEM[37147] + MEM[37256];
assign MEM[43507] = MEM[37149] + MEM[37248];
assign MEM[43508] = MEM[37152] + MEM[37210];
assign MEM[43509] = MEM[37153] + MEM[37306];
assign MEM[43510] = MEM[37154] + MEM[37296];
assign MEM[43511] = MEM[37156] + MEM[37190];
assign MEM[43512] = MEM[37158] + MEM[37203];
assign MEM[43513] = MEM[37160] + MEM[37218];
assign MEM[43514] = MEM[37161] + MEM[37169];
assign MEM[43515] = MEM[37163] + MEM[37199];
assign MEM[43516] = MEM[37164] + MEM[37187];
assign MEM[43517] = MEM[37166] + MEM[37170];
assign MEM[43518] = MEM[37167] + MEM[37192];
assign MEM[43519] = MEM[37168] + MEM[37216];
assign MEM[43520] = MEM[37172] + MEM[37249];
assign MEM[43521] = MEM[37174] + MEM[37259];
assign MEM[43522] = MEM[37175] + MEM[37193];
assign MEM[43523] = MEM[37176] + MEM[37271];
assign MEM[43524] = MEM[37177] + MEM[37207];
assign MEM[43525] = MEM[37178] + MEM[37253];
assign MEM[43526] = MEM[37180] + MEM[37228];
assign MEM[43527] = MEM[37181] + MEM[37208];
assign MEM[43528] = MEM[37183] + MEM[37220];
assign MEM[43529] = MEM[37185] + MEM[37197];
assign MEM[43530] = MEM[37186] + MEM[37202];
assign MEM[43531] = MEM[37194] + MEM[37233];
assign MEM[43532] = MEM[37195] + MEM[37239];
assign MEM[43533] = MEM[37196] + MEM[37321];
assign MEM[43534] = MEM[37200] + MEM[37235];
assign MEM[43535] = MEM[37204] + MEM[37237];
assign MEM[43536] = MEM[37205] + MEM[37298];
assign MEM[43537] = MEM[37206] + MEM[37275];
assign MEM[43538] = MEM[37209] + MEM[37226];
assign MEM[43539] = MEM[37212] + MEM[37286];
assign MEM[43540] = MEM[37213] + MEM[37304];
assign MEM[43541] = MEM[37215] + MEM[37345];
assign MEM[43542] = MEM[37217] + MEM[37245];
assign MEM[43543] = MEM[37219] + MEM[37308];
assign MEM[43544] = MEM[37221] + MEM[37299];
assign MEM[43545] = MEM[37222] + MEM[37391];
assign MEM[43546] = MEM[37224] + MEM[37243];
assign MEM[43547] = MEM[37225] + MEM[37287];
assign MEM[43548] = MEM[37229] + MEM[37288];
assign MEM[43549] = MEM[37230] + MEM[37247];
assign MEM[43550] = MEM[37231] + MEM[37336];
assign MEM[43551] = MEM[37234] + MEM[37369];
assign MEM[43552] = MEM[37236] + MEM[37278];
assign MEM[43553] = MEM[37240] + MEM[37269];
assign MEM[43554] = MEM[37244] + MEM[37370];
assign MEM[43555] = MEM[37250] + MEM[37397];
assign MEM[43556] = MEM[37251] + MEM[37291];
assign MEM[43557] = MEM[37252] + MEM[37284];
assign MEM[43558] = MEM[37254] + MEM[37385];
assign MEM[43559] = MEM[37255] + MEM[37297];
assign MEM[43560] = MEM[37258] + MEM[37407];
assign MEM[43561] = MEM[37260] + MEM[37280];
assign MEM[43562] = MEM[37261] + MEM[37316];
assign MEM[43563] = MEM[37262] + MEM[37281];
assign MEM[43564] = MEM[37263] + MEM[37422];
assign MEM[43565] = MEM[37264] + MEM[37386];
assign MEM[43566] = MEM[37265] + MEM[37313];
assign MEM[43567] = MEM[37266] + MEM[37320];
assign MEM[43568] = MEM[37267] + MEM[37390];
assign MEM[43569] = MEM[37268] + MEM[37373];
assign MEM[43570] = MEM[37270] + MEM[37358];
assign MEM[43571] = MEM[37272] + MEM[37305];
assign MEM[43572] = MEM[37273] + MEM[37301];
assign MEM[43573] = MEM[37274] + MEM[37311];
assign MEM[43574] = MEM[37276] + MEM[37339];
assign MEM[43575] = MEM[37277] + MEM[37327];
assign MEM[43576] = MEM[37279] + MEM[37295];
assign MEM[43577] = MEM[37282] + MEM[37335];
assign MEM[43578] = MEM[37283] + MEM[37314];
assign MEM[43579] = MEM[37285] + MEM[37303];
assign MEM[43580] = MEM[37290] + MEM[37302];
assign MEM[43581] = MEM[37292] + MEM[37319];
assign MEM[43582] = MEM[37293] + MEM[37315];
assign MEM[43583] = MEM[37294] + MEM[37387];
assign MEM[43584] = MEM[37300] + MEM[37353];
assign MEM[43585] = MEM[37307] + MEM[37328];
assign MEM[43586] = MEM[37309] + MEM[37324];
assign MEM[43587] = MEM[37310] + MEM[37444];
assign MEM[43588] = MEM[37312] + MEM[37406];
assign MEM[43589] = MEM[37317] + MEM[37522];
assign MEM[43590] = MEM[37318] + MEM[37338];
assign MEM[43591] = MEM[37322] + MEM[37383];
assign MEM[43592] = MEM[37323] + MEM[37416];
assign MEM[43593] = MEM[37325] + MEM[37366];
assign MEM[43594] = MEM[37329] + MEM[37372];
assign MEM[43595] = MEM[37330] + MEM[37481];
assign MEM[43596] = MEM[37331] + MEM[37360];
assign MEM[43597] = MEM[37332] + MEM[37346];
assign MEM[43598] = MEM[37333] + MEM[37356];
assign MEM[43599] = MEM[37334] + MEM[37409];
assign MEM[43600] = MEM[37337] + MEM[37418];
assign MEM[43601] = MEM[37340] + MEM[37414];
assign MEM[43602] = MEM[37341] + MEM[37446];
assign MEM[43603] = MEM[37342] + MEM[37393];
assign MEM[43604] = MEM[37343] + MEM[37455];
assign MEM[43605] = MEM[37344] + MEM[37412];
assign MEM[43606] = MEM[37347] + MEM[37349];
assign MEM[43607] = MEM[37348] + MEM[37381];
assign MEM[43608] = MEM[37350] + MEM[37392];
assign MEM[43609] = MEM[37351] + MEM[37505];
assign MEM[43610] = MEM[37352] + MEM[37380];
assign MEM[43611] = MEM[37354] + MEM[37364];
assign MEM[43612] = MEM[37355] + MEM[37362];
assign MEM[43613] = MEM[37357] + MEM[37430];
assign MEM[43614] = MEM[37359] + MEM[37396];
assign MEM[43615] = MEM[37361] + MEM[37411];
assign MEM[43616] = MEM[37363] + MEM[37403];
assign MEM[43617] = MEM[37365] + MEM[37436];
assign MEM[43618] = MEM[37367] + MEM[37402];
assign MEM[43619] = MEM[37368] + MEM[37434];
assign MEM[43620] = MEM[37371] + MEM[37472];
assign MEM[43621] = MEM[37374] + MEM[37419];
assign MEM[43622] = MEM[37375] + MEM[37442];
assign MEM[43623] = MEM[37376] + MEM[37423];
assign MEM[43624] = MEM[37377] + MEM[37382];
assign MEM[43625] = MEM[37378] + MEM[37476];
assign MEM[43626] = MEM[37379] + MEM[37469];
assign MEM[43627] = MEM[37384] + MEM[37432];
assign MEM[43628] = MEM[37388] + MEM[37428];
assign MEM[43629] = MEM[37389] + MEM[37433];
assign MEM[43630] = MEM[37394] + MEM[37401];
assign MEM[43631] = MEM[37395] + MEM[37415];
assign MEM[43632] = MEM[37398] + MEM[37467];
assign MEM[43633] = MEM[37399] + MEM[37536];
assign MEM[43634] = MEM[37400] + MEM[37462];
assign MEM[43635] = MEM[37404] + MEM[37486];
assign MEM[43636] = MEM[37405] + MEM[37484];
assign MEM[43637] = MEM[37408] + MEM[37463];
assign MEM[43638] = MEM[37410] + MEM[37453];
assign MEM[43639] = MEM[37413] + MEM[37452];
assign MEM[43640] = MEM[37417] + MEM[37445];
assign MEM[43641] = MEM[37420] + MEM[37431];
assign MEM[43642] = MEM[37421] + MEM[37479];
assign MEM[43643] = MEM[37424] + MEM[37567];
assign MEM[43644] = MEM[37425] + MEM[37451];
assign MEM[43645] = MEM[37426] + MEM[37518];
assign MEM[43646] = MEM[37427] + MEM[37509];
assign MEM[43647] = MEM[37429] + MEM[37517];
assign MEM[43648] = MEM[37435] + MEM[37470];
assign MEM[43649] = MEM[37437] + MEM[37573];
assign MEM[43650] = MEM[37438] + MEM[37483];
assign MEM[43651] = MEM[37439] + MEM[37540];
assign MEM[43652] = MEM[37440] + MEM[37526];
assign MEM[43653] = MEM[37441] + MEM[37495];
assign MEM[43654] = MEM[37443] + MEM[37533];
assign MEM[43655] = MEM[37447] + MEM[37569];
assign MEM[43656] = MEM[37448] + MEM[37530];
assign MEM[43657] = MEM[37449] + MEM[37497];
assign MEM[43658] = MEM[37450] + MEM[37514];
assign MEM[43659] = MEM[37454] + MEM[37538];
assign MEM[43660] = MEM[37456] + MEM[37501];
assign MEM[43661] = MEM[37457] + MEM[37494];
assign MEM[43662] = MEM[37458] + MEM[37465];
assign MEM[43663] = MEM[37459] + MEM[37549];
assign MEM[43664] = MEM[37460] + MEM[37488];
assign MEM[43665] = MEM[37461] + MEM[37576];
assign MEM[43666] = MEM[37464] + MEM[37524];
assign MEM[43667] = MEM[37466] + MEM[37512];
assign MEM[43668] = MEM[37468] + MEM[37508];
assign MEM[43669] = MEM[37471] + MEM[37565];
assign MEM[43670] = MEM[37473] + MEM[37493];
assign MEM[43671] = MEM[37474] + MEM[37582];
assign MEM[43672] = MEM[37475] + MEM[37527];
assign MEM[43673] = MEM[37477] + MEM[37489];
assign MEM[43674] = MEM[37478] + MEM[37492];
assign MEM[43675] = MEM[37480] + MEM[37571];
assign MEM[43676] = MEM[37482] + MEM[37546];
assign MEM[43677] = MEM[37485] + MEM[37541];
assign MEM[43678] = MEM[37487] + MEM[37516];
assign MEM[43679] = MEM[37490] + MEM[37507];
assign MEM[43680] = MEM[37491] + MEM[37531];
assign MEM[43681] = MEM[37496] + MEM[37523];
assign MEM[43682] = MEM[37498] + MEM[37578];
assign MEM[43683] = MEM[37499] + MEM[37638];
assign MEM[43684] = MEM[37500] + MEM[37520];
assign MEM[43685] = MEM[37502] + MEM[37606];
assign MEM[43686] = MEM[37503] + MEM[37589];
assign MEM[43687] = MEM[37504] + MEM[37684];
assign MEM[43688] = MEM[37506] + MEM[37521];
assign MEM[43689] = MEM[37510] + MEM[37563];
assign MEM[43690] = MEM[37511] + MEM[37598];
assign MEM[43691] = MEM[37513] + MEM[37545];
assign MEM[43692] = MEM[37515] + MEM[37566];
assign MEM[43693] = MEM[37519] + MEM[37622];
assign MEM[43694] = MEM[37525] + MEM[37602];
assign MEM[43695] = MEM[37528] + MEM[37644];
assign MEM[43696] = MEM[37529] + MEM[37543];
assign MEM[43697] = MEM[37532] + MEM[37605];
assign MEM[43698] = MEM[37534] + MEM[37556];
assign MEM[43699] = MEM[37535] + MEM[37619];
assign MEM[43700] = MEM[37537] + MEM[37610];
assign MEM[43701] = MEM[37539] + MEM[37681];
assign MEM[43702] = MEM[37542] + MEM[37561];
assign MEM[43703] = MEM[37544] + MEM[37557];
assign MEM[43704] = MEM[37547] + MEM[37662];
assign MEM[43705] = MEM[37548] + MEM[37593];
assign MEM[43706] = MEM[37550] + MEM[37596];
assign MEM[43707] = MEM[37551] + MEM[37600];
assign MEM[43708] = MEM[37552] + MEM[37625];
assign MEM[43709] = MEM[37553] + MEM[37654];
assign MEM[43710] = MEM[37554] + MEM[37590];
assign MEM[43711] = MEM[37555] + MEM[37591];
assign MEM[43712] = MEM[37558] + MEM[37620];
assign MEM[43713] = MEM[37559] + MEM[37617];
assign MEM[43714] = MEM[37560] + MEM[37583];
assign MEM[43715] = MEM[37562] + MEM[37597];
assign MEM[43716] = MEM[37564] + MEM[37584];
assign MEM[43717] = MEM[37568] + MEM[37608];
assign MEM[43718] = MEM[37570] + MEM[37672];
assign MEM[43719] = MEM[37572] + MEM[37604];
assign MEM[43720] = MEM[37574] + MEM[37643];
assign MEM[43721] = MEM[37575] + MEM[37666];
assign MEM[43722] = MEM[37577] + MEM[37674];
assign MEM[43723] = MEM[37579] + MEM[37718];
assign MEM[43724] = MEM[37580] + MEM[37613];
assign MEM[43725] = MEM[37581] + MEM[37664];
assign MEM[43726] = MEM[37585] + MEM[37685];
assign MEM[43727] = MEM[37586] + MEM[37642];
assign MEM[43728] = MEM[37587] + MEM[37663];
assign MEM[43729] = MEM[37588] + MEM[37603];
assign MEM[43730] = MEM[37592] + MEM[37677];
assign MEM[43731] = MEM[37594] + MEM[37631];
assign MEM[43732] = MEM[37595] + MEM[37687];
assign MEM[43733] = MEM[37599] + MEM[37669];
assign MEM[43734] = MEM[37601] + MEM[37648];
assign MEM[43735] = MEM[37607] + MEM[37826];
assign MEM[43736] = MEM[37609] + MEM[37975];
assign MEM[43737] = MEM[37611] + MEM[37657];
assign MEM[43738] = MEM[37612] + MEM[37660];
assign MEM[43739] = MEM[37614] + MEM[37700];
assign MEM[43740] = MEM[37615] + MEM[37628];
assign MEM[43741] = MEM[37616] + MEM[37692];
assign MEM[43742] = MEM[37618] + MEM[37713];
assign MEM[43743] = MEM[37621] + MEM[37704];
assign MEM[43744] = MEM[37623] + MEM[37731];
assign MEM[43745] = MEM[37624] + MEM[37693];
assign MEM[43746] = MEM[37626] + MEM[37719];
assign MEM[43747] = MEM[37627] + MEM[37679];
assign MEM[43748] = MEM[37629] + MEM[37640];
assign MEM[43749] = MEM[37630] + MEM[37652];
assign MEM[43750] = MEM[37632] + MEM[37747];
assign MEM[43751] = MEM[37633] + MEM[37678];
assign MEM[43752] = MEM[37634] + MEM[37686];
assign MEM[43753] = MEM[37635] + MEM[37667];
assign MEM[43754] = MEM[37636] + MEM[37701];
assign MEM[43755] = MEM[37637] + MEM[37734];
assign MEM[43756] = MEM[37639] + MEM[37653];
assign MEM[43757] = MEM[37641] + MEM[37698];
assign MEM[43758] = MEM[37645] + MEM[37697];
assign MEM[43759] = MEM[37646] + MEM[37694];
assign MEM[43760] = MEM[37647] + MEM[37661];
assign MEM[43761] = MEM[37649] + MEM[37720];
assign MEM[43762] = MEM[37650] + MEM[37671];
assign MEM[43763] = MEM[37651] + MEM[37696];
assign MEM[43764] = MEM[37655] + MEM[37715];
assign MEM[43765] = MEM[37656] + MEM[37785];
assign MEM[43766] = MEM[37658] + MEM[37709];
assign MEM[43767] = MEM[37659] + MEM[37675];
assign MEM[43768] = MEM[37665] + MEM[37844];
assign MEM[43769] = MEM[37668] + MEM[37723];
assign MEM[43770] = MEM[37670] + MEM[37764];
assign MEM[43771] = MEM[37673] + MEM[37707];
assign MEM[43772] = MEM[37676] + MEM[37732];
assign MEM[43773] = MEM[37680] + MEM[37724];
assign MEM[43774] = MEM[37682] + MEM[37827];
assign MEM[43775] = MEM[37683] + MEM[37691];
assign MEM[43776] = MEM[37688] + MEM[37752];
assign MEM[43777] = MEM[37689] + MEM[37710];
assign MEM[43778] = MEM[37690] + MEM[37725];
assign MEM[43779] = MEM[37695] + MEM[37781];
assign MEM[43780] = MEM[37699] + MEM[37750];
assign MEM[43781] = MEM[37702] + MEM[37728];
assign MEM[43782] = MEM[37703] + MEM[37882];
assign MEM[43783] = MEM[37705] + MEM[37748];
assign MEM[43784] = MEM[37706] + MEM[37765];
assign MEM[43785] = MEM[37708] + MEM[37760];
assign MEM[43786] = MEM[37711] + MEM[37761];
assign MEM[43787] = MEM[37712] + MEM[37758];
assign MEM[43788] = MEM[37714] + MEM[37816];
assign MEM[43789] = MEM[37716] + MEM[37756];
assign MEM[43790] = MEM[37717] + MEM[37763];
assign MEM[43791] = MEM[37721] + MEM[37782];
assign MEM[43792] = MEM[37722] + MEM[37757];
assign MEM[43793] = MEM[37726] + MEM[37776];
assign MEM[43794] = MEM[37727] + MEM[37770];
assign MEM[43795] = MEM[37729] + MEM[37766];
assign MEM[43796] = MEM[37730] + MEM[37783];
assign MEM[43797] = MEM[37733] + MEM[37762];
assign MEM[43798] = MEM[37735] + MEM[37853];
assign MEM[43799] = MEM[37736] + MEM[37804];
assign MEM[43800] = MEM[37737] + MEM[37769];
assign MEM[43801] = MEM[37738] + MEM[37778];
assign MEM[43802] = MEM[37739] + MEM[37772];
assign MEM[43803] = MEM[37740] + MEM[37822];
assign MEM[43804] = MEM[37741] + MEM[37796];
assign MEM[43805] = MEM[37742] + MEM[37802];
assign MEM[43806] = MEM[37743] + MEM[37848];
assign MEM[43807] = MEM[37744] + MEM[37786];
assign MEM[43808] = MEM[37745] + MEM[37795];
assign MEM[43809] = MEM[37746] + MEM[37800];
assign MEM[43810] = MEM[37749] + MEM[37771];
assign MEM[43811] = MEM[37751] + MEM[37851];
assign MEM[43812] = MEM[37753] + MEM[37830];
assign MEM[43813] = MEM[37754] + MEM[37774];
assign MEM[43814] = MEM[37755] + MEM[37798];
assign MEM[43815] = MEM[37759] + MEM[37865];
assign MEM[43816] = MEM[37767] + MEM[37897];
assign MEM[43817] = MEM[37768] + MEM[37817];
assign MEM[43818] = MEM[37773] + MEM[37835];
assign MEM[43819] = MEM[37775] + MEM[37818];
assign MEM[43820] = MEM[37777] + MEM[37916];
assign MEM[43821] = MEM[37779] + MEM[37863];
assign MEM[43822] = MEM[37780] + MEM[37793];
assign MEM[43823] = MEM[37784] + MEM[37808];
assign MEM[43824] = MEM[37787] + MEM[37860];
assign MEM[43825] = MEM[37788] + MEM[37831];
assign MEM[43826] = MEM[37789] + MEM[37824];
assign MEM[43827] = MEM[37790] + MEM[37942];
assign MEM[43828] = MEM[37791] + MEM[37854];
assign MEM[43829] = MEM[37792] + MEM[37820];
assign MEM[43830] = MEM[37794] + MEM[37950];
assign MEM[43831] = MEM[37797] + MEM[37862];
assign MEM[43832] = MEM[37799] + MEM[37811];
assign MEM[43833] = MEM[37801] + MEM[38032];
assign MEM[43834] = MEM[37803] + MEM[37849];
assign MEM[43835] = MEM[37805] + MEM[37834];
assign MEM[43836] = MEM[37806] + MEM[37912];
assign MEM[43837] = MEM[37807] + MEM[37869];
assign MEM[43838] = MEM[37809] + MEM[37825];
assign MEM[43839] = MEM[37810] + MEM[37928];
assign MEM[43840] = MEM[37812] + MEM[37858];
assign MEM[43841] = MEM[37813] + MEM[37935];
assign MEM[43842] = MEM[37814] + MEM[37871];
assign MEM[43843] = MEM[37815] + MEM[37955];
assign MEM[43844] = MEM[37819] + MEM[37859];
assign MEM[43845] = MEM[37821] + MEM[37976];
assign MEM[43846] = MEM[37823] + MEM[37881];
assign MEM[43847] = MEM[37828] + MEM[38005];
assign MEM[43848] = MEM[37829] + MEM[37884];
assign MEM[43849] = MEM[37832] + MEM[37899];
assign MEM[43850] = MEM[37833] + MEM[37878];
assign MEM[43851] = MEM[37836] + MEM[37988];
assign MEM[43852] = MEM[37837] + MEM[37887];
assign MEM[43853] = MEM[37838] + MEM[37900];
assign MEM[43854] = MEM[37839] + MEM[37876];
assign MEM[43855] = MEM[37840] + MEM[37879];
assign MEM[43856] = MEM[37841] + MEM[37872];
assign MEM[43857] = MEM[37842] + MEM[37906];
assign MEM[43858] = MEM[37843] + MEM[37902];
assign MEM[43859] = MEM[37845] + MEM[37885];
assign MEM[43860] = MEM[37846] + MEM[37901];
assign MEM[43861] = MEM[37847] + MEM[37964];
assign MEM[43862] = MEM[37850] + MEM[37864];
assign MEM[43863] = MEM[37852] + MEM[37948];
assign MEM[43864] = MEM[37855] + MEM[37880];
assign MEM[43865] = MEM[37856] + MEM[37875];
assign MEM[43866] = MEM[37857] + MEM[37891];
assign MEM[43867] = MEM[37861] + MEM[38081];
assign MEM[43868] = MEM[37866] + MEM[37893];
assign MEM[43869] = MEM[37867] + MEM[37914];
assign MEM[43870] = MEM[37868] + MEM[37883];
assign MEM[43871] = MEM[37870] + MEM[37915];
assign MEM[43872] = MEM[37873] + MEM[37965];
assign MEM[43873] = MEM[37874] + MEM[37922];
assign MEM[43874] = MEM[37877] + MEM[37984];
assign MEM[43875] = MEM[37886] + MEM[37911];
assign MEM[43876] = MEM[37888] + MEM[38038];
assign MEM[43877] = MEM[37889] + MEM[37968];
assign MEM[43878] = MEM[37890] + MEM[38001];
assign MEM[43879] = MEM[37892] + MEM[37904];
assign MEM[43880] = MEM[37894] + MEM[37923];
assign MEM[43881] = MEM[37895] + MEM[38022];
assign MEM[43882] = MEM[37896] + MEM[37995];
assign MEM[43883] = MEM[37898] + MEM[38000];
assign MEM[43884] = MEM[37903] + MEM[37989];
assign MEM[43885] = MEM[37905] + MEM[38006];
assign MEM[43886] = MEM[37907] + MEM[37993];
assign MEM[43887] = MEM[37908] + MEM[37971];
assign MEM[43888] = MEM[37909] + MEM[37986];
assign MEM[43889] = MEM[37910] + MEM[37951];
assign MEM[43890] = MEM[37913] + MEM[37941];
assign MEM[43891] = MEM[37917] + MEM[37947];
assign MEM[43892] = MEM[37918] + MEM[37946];
assign MEM[43893] = MEM[37919] + MEM[37952];
assign MEM[43894] = MEM[37920] + MEM[37956];
assign MEM[43895] = MEM[37921] + MEM[37926];
assign MEM[43896] = MEM[37924] + MEM[37930];
assign MEM[43897] = MEM[37925] + MEM[38017];
assign MEM[43898] = MEM[37927] + MEM[37962];
assign MEM[43899] = MEM[37929] + MEM[37958];
assign MEM[43900] = MEM[37931] + MEM[37985];
assign MEM[43901] = MEM[37932] + MEM[37982];
assign MEM[43902] = MEM[37933] + MEM[37949];
assign MEM[43903] = MEM[37934] + MEM[37957];
assign MEM[43904] = MEM[37936] + MEM[38039];
assign MEM[43905] = MEM[37937] + MEM[37966];
assign MEM[43906] = MEM[37938] + MEM[38035];
assign MEM[43907] = MEM[37939] + MEM[37960];
assign MEM[43908] = MEM[37940] + MEM[37959];
assign MEM[43909] = MEM[37943] + MEM[38082];
assign MEM[43910] = MEM[37944] + MEM[38030];
assign MEM[43911] = MEM[37945] + MEM[38024];
assign MEM[43912] = MEM[37953] + MEM[38031];
assign MEM[43913] = MEM[37954] + MEM[38011];
assign MEM[43914] = MEM[37961] + MEM[37997];
assign MEM[43915] = MEM[37963] + MEM[37983];
assign MEM[43916] = MEM[37967] + MEM[38037];
assign MEM[43917] = MEM[37969] + MEM[38028];
assign MEM[43918] = MEM[37970] + MEM[38004];
assign MEM[43919] = MEM[37972] + MEM[38019];
assign MEM[43920] = MEM[37973] + MEM[38044];
assign MEM[43921] = MEM[37974] + MEM[38051];
assign MEM[43922] = MEM[37977] + MEM[38047];
assign MEM[43923] = MEM[37978] + MEM[38118];
assign MEM[43924] = MEM[37979] + MEM[38021];
assign MEM[43925] = MEM[37980] + MEM[38066];
assign MEM[43926] = MEM[37981] + MEM[38069];
assign MEM[43927] = MEM[37987] + MEM[38033];
assign MEM[43928] = MEM[37990] + MEM[38020];
assign MEM[43929] = MEM[37991] + MEM[38113];
assign MEM[43930] = MEM[37992] + MEM[38109];
assign MEM[43931] = MEM[37994] + MEM[38115];
assign MEM[43932] = MEM[37996] + MEM[38104];
assign MEM[43933] = MEM[37998] + MEM[38013];
assign MEM[43934] = MEM[37999] + MEM[38034];
assign MEM[43935] = MEM[38002] + MEM[38106];
assign MEM[43936] = MEM[38003] + MEM[38043];
assign MEM[43937] = MEM[38007] + MEM[38015];
assign MEM[43938] = MEM[38008] + MEM[38056];
assign MEM[43939] = MEM[38009] + MEM[38079];
assign MEM[43940] = MEM[38010] + MEM[38027];
assign MEM[43941] = MEM[38012] + MEM[38067];
assign MEM[43942] = MEM[38014] + MEM[38132];
assign MEM[43943] = MEM[38016] + MEM[38042];
assign MEM[43944] = MEM[38018] + MEM[38046];
assign MEM[43945] = MEM[38023] + MEM[38119];
assign MEM[43946] = MEM[38025] + MEM[38126];
assign MEM[43947] = MEM[38026] + MEM[38101];
assign MEM[43948] = MEM[38029] + MEM[38108];
assign MEM[43949] = MEM[38036] + MEM[38052];
assign MEM[43950] = MEM[38040] + MEM[38135];
assign MEM[43951] = MEM[38041] + MEM[38159];
assign MEM[43952] = MEM[38045] + MEM[38049];
assign MEM[43953] = MEM[38048] + MEM[38080];
assign MEM[43954] = MEM[38050] + MEM[38092];
assign MEM[43955] = MEM[38053] + MEM[38160];
assign MEM[43956] = MEM[38054] + MEM[38073];
assign MEM[43957] = MEM[38055] + MEM[38099];
assign MEM[43958] = MEM[38057] + MEM[38068];
assign MEM[43959] = MEM[38058] + MEM[38071];
assign MEM[43960] = MEM[38059] + MEM[38100];
assign MEM[43961] = MEM[38060] + MEM[38093];
assign MEM[43962] = MEM[38061] + MEM[38077];
assign MEM[43963] = MEM[38062] + MEM[38179];
assign MEM[43964] = MEM[38063] + MEM[38112];
assign MEM[43965] = MEM[38064] + MEM[38149];
assign MEM[43966] = MEM[38065] + MEM[38107];
assign MEM[43967] = MEM[38070] + MEM[38105];
assign MEM[43968] = MEM[38072] + MEM[38154];
assign MEM[43969] = MEM[38074] + MEM[38166];
assign MEM[43970] = MEM[38075] + MEM[38251];
assign MEM[43971] = MEM[38076] + MEM[38136];
assign MEM[43972] = MEM[38078] + MEM[38134];
assign MEM[43973] = MEM[38083] + MEM[38095];
assign MEM[43974] = MEM[38084] + MEM[38117];
assign MEM[43975] = MEM[38085] + MEM[38125];
assign MEM[43976] = MEM[38086] + MEM[38172];
assign MEM[43977] = MEM[38087] + MEM[38196];
assign MEM[43978] = MEM[38088] + MEM[38194];
assign MEM[43979] = MEM[38089] + MEM[38204];
assign MEM[43980] = MEM[38090] + MEM[38140];
assign MEM[43981] = MEM[38091] + MEM[38153];
assign MEM[43982] = MEM[38094] + MEM[38175];
assign MEM[43983] = MEM[38096] + MEM[38222];
assign MEM[43984] = MEM[38097] + MEM[38111];
assign MEM[43985] = MEM[38098] + MEM[38152];
assign MEM[43986] = MEM[38102] + MEM[38215];
assign MEM[43987] = MEM[38103] + MEM[38190];
assign MEM[43988] = MEM[38110] + MEM[38203];
assign MEM[43989] = MEM[38114] + MEM[38151];
assign MEM[43990] = MEM[38116] + MEM[38148];
assign MEM[43991] = MEM[38120] + MEM[38147];
assign MEM[43992] = MEM[38121] + MEM[38164];
assign MEM[43993] = MEM[38122] + MEM[38169];
assign MEM[43994] = MEM[38123] + MEM[38176];
assign MEM[43995] = MEM[38124] + MEM[38209];
assign MEM[43996] = MEM[38127] + MEM[38163];
assign MEM[43997] = MEM[38128] + MEM[38185];
assign MEM[43998] = MEM[38129] + MEM[38188];
assign MEM[43999] = MEM[38130] + MEM[38177];
assign MEM[44000] = MEM[38131] + MEM[38146];
assign MEM[44001] = MEM[38133] + MEM[38174];
assign MEM[44002] = MEM[38137] + MEM[38221];
assign MEM[44003] = MEM[38138] + MEM[38212];
assign MEM[44004] = MEM[38139] + MEM[38173];
assign MEM[44005] = MEM[38141] + MEM[38220];
assign MEM[44006] = MEM[38142] + MEM[38202];
assign MEM[44007] = MEM[38143] + MEM[38187];
assign MEM[44008] = MEM[38144] + MEM[38223];
assign MEM[44009] = MEM[38145] + MEM[38218];
assign MEM[44010] = MEM[38150] + MEM[38156];
assign MEM[44011] = MEM[38155] + MEM[38168];
assign MEM[44012] = MEM[38157] + MEM[38265];
assign MEM[44013] = MEM[38158] + MEM[38191];
assign MEM[44014] = MEM[38161] + MEM[38264];
assign MEM[44015] = MEM[38162] + MEM[38226];
assign MEM[44016] = MEM[38165] + MEM[38259];
assign MEM[44017] = MEM[38167] + MEM[38214];
assign MEM[44018] = MEM[38170] + MEM[38276];
assign MEM[44019] = MEM[38171] + MEM[38205];
assign MEM[44020] = MEM[38178] + MEM[38183];
assign MEM[44021] = MEM[38180] + MEM[38355];
assign MEM[44022] = MEM[38181] + MEM[38238];
assign MEM[44023] = MEM[38182] + MEM[38245];
assign MEM[44024] = MEM[38184] + MEM[38239];
assign MEM[44025] = MEM[38186] + MEM[38288];
assign MEM[44026] = MEM[38189] + MEM[38320];
assign MEM[44027] = MEM[38192] + MEM[38309];
assign MEM[44028] = MEM[38193] + MEM[38213];
assign MEM[44029] = MEM[38195] + MEM[38208];
assign MEM[44030] = MEM[38197] + MEM[38252];
assign MEM[44031] = MEM[38198] + MEM[38224];
assign MEM[44032] = MEM[38199] + MEM[38227];
assign MEM[44033] = MEM[38200] + MEM[38302];
assign MEM[44034] = MEM[38201] + MEM[38237];
assign MEM[44035] = MEM[38206] + MEM[38275];
assign MEM[44036] = MEM[38207] + MEM[38247];
assign MEM[44037] = MEM[38210] + MEM[38271];
assign MEM[44038] = MEM[38211] + MEM[38232];
assign MEM[44039] = MEM[38216] + MEM[38249];
assign MEM[44040] = MEM[38217] + MEM[38304];
assign MEM[44041] = MEM[38219] + MEM[38329];
assign MEM[44042] = MEM[38225] + MEM[38233];
assign MEM[44043] = MEM[38228] + MEM[38373];
assign MEM[44044] = MEM[38229] + MEM[38256];
assign MEM[44045] = MEM[38230] + MEM[38319];
assign MEM[44046] = MEM[38231] + MEM[38250];
assign MEM[44047] = MEM[38234] + MEM[38299];
assign MEM[44048] = MEM[38235] + MEM[38522];
assign MEM[44049] = MEM[38236] + MEM[38405];
assign MEM[44050] = MEM[38240] + MEM[38316];
assign MEM[44051] = MEM[38241] + MEM[38325];
assign MEM[44052] = MEM[38242] + MEM[38310];
assign MEM[44053] = MEM[38243] + MEM[38311];
assign MEM[44054] = MEM[38244] + MEM[38286];
assign MEM[44055] = MEM[38246] + MEM[38261];
assign MEM[44056] = MEM[38248] + MEM[38305];
assign MEM[44057] = MEM[38253] + MEM[38287];
assign MEM[44058] = MEM[38254] + MEM[38269];
assign MEM[44059] = MEM[38255] + MEM[38343];
assign MEM[44060] = MEM[38257] + MEM[38348];
assign MEM[44061] = MEM[38258] + MEM[38317];
assign MEM[44062] = MEM[38260] + MEM[38301];
assign MEM[44063] = MEM[38262] + MEM[38308];
assign MEM[44064] = MEM[38263] + MEM[38389];
assign MEM[44065] = MEM[38266] + MEM[38367];
assign MEM[44066] = MEM[38267] + MEM[38298];
assign MEM[44067] = MEM[38268] + MEM[38291];
assign MEM[44068] = MEM[38270] + MEM[38292];
assign MEM[44069] = MEM[38272] + MEM[38378];
assign MEM[44070] = MEM[38273] + MEM[38323];
assign MEM[44071] = MEM[38274] + MEM[38341];
assign MEM[44072] = MEM[38277] + MEM[38339];
assign MEM[44073] = MEM[38278] + MEM[38377];
assign MEM[44074] = MEM[38279] + MEM[38331];
assign MEM[44075] = MEM[38280] + MEM[38318];
assign MEM[44076] = MEM[38281] + MEM[38321];
assign MEM[44077] = MEM[38282] + MEM[38296];
assign MEM[44078] = MEM[38283] + MEM[38297];
assign MEM[44079] = MEM[38284] + MEM[38315];
assign MEM[44080] = MEM[38285] + MEM[38324];
assign MEM[44081] = MEM[38289] + MEM[38431];
assign MEM[44082] = MEM[38290] + MEM[38399];
assign MEM[44083] = MEM[38293] + MEM[38362];
assign MEM[44084] = MEM[38294] + MEM[38411];
assign MEM[44085] = MEM[38295] + MEM[38372];
assign MEM[44086] = MEM[38300] + MEM[38387];
assign MEM[44087] = MEM[38303] + MEM[38393];
assign MEM[44088] = MEM[38306] + MEM[38337];
assign MEM[44089] = MEM[38307] + MEM[38379];
assign MEM[44090] = MEM[38312] + MEM[38342];
assign MEM[44091] = MEM[38313] + MEM[38335];
assign MEM[44092] = MEM[38314] + MEM[38385];
assign MEM[44093] = MEM[38322] + MEM[38388];
assign MEM[44094] = MEM[38326] + MEM[38427];
assign MEM[44095] = MEM[38327] + MEM[38382];
assign MEM[44096] = MEM[38328] + MEM[38419];
assign MEM[44097] = MEM[38330] + MEM[38361];
assign MEM[44098] = MEM[38332] + MEM[38420];
assign MEM[44099] = MEM[38333] + MEM[38357];
assign MEM[44100] = MEM[38334] + MEM[38457];
assign MEM[44101] = MEM[38336] + MEM[38349];
assign MEM[44102] = MEM[38338] + MEM[38368];
assign MEM[44103] = MEM[38340] + MEM[38365];
assign MEM[44104] = MEM[38344] + MEM[38446];
assign MEM[44105] = MEM[38345] + MEM[38364];
assign MEM[44106] = MEM[38346] + MEM[38423];
assign MEM[44107] = MEM[38347] + MEM[38408];
assign MEM[44108] = MEM[38350] + MEM[38406];
assign MEM[44109] = MEM[38351] + MEM[38394];
assign MEM[44110] = MEM[38352] + MEM[38402];
assign MEM[44111] = MEM[38353] + MEM[38413];
assign MEM[44112] = MEM[38354] + MEM[38386];
assign MEM[44113] = MEM[38356] + MEM[38384];
assign MEM[44114] = MEM[38358] + MEM[38418];
assign MEM[44115] = MEM[38359] + MEM[38375];
assign MEM[44116] = MEM[38360] + MEM[38398];
assign MEM[44117] = MEM[38363] + MEM[38443];
assign MEM[44118] = MEM[38366] + MEM[38403];
assign MEM[44119] = MEM[38369] + MEM[38416];
assign MEM[44120] = MEM[38370] + MEM[38517];
assign MEM[44121] = MEM[38371] + MEM[38435];
assign MEM[44122] = MEM[38374] + MEM[38395];
assign MEM[44123] = MEM[38376] + MEM[38448];
assign MEM[44124] = MEM[38380] + MEM[38415];
assign MEM[44125] = MEM[38381] + MEM[38483];
assign MEM[44126] = MEM[38383] + MEM[38414];
assign MEM[44127] = MEM[38390] + MEM[38498];
assign MEM[44128] = MEM[38391] + MEM[38409];
assign MEM[44129] = MEM[38392] + MEM[38467];
assign MEM[44130] = MEM[38396] + MEM[38429];
assign MEM[44131] = MEM[38397] + MEM[38468];
assign MEM[44132] = MEM[38400] + MEM[38452];
assign MEM[44133] = MEM[38401] + MEM[38473];
assign MEM[44134] = MEM[38404] + MEM[38426];
assign MEM[44135] = MEM[38407] + MEM[38543];
assign MEM[44136] = MEM[38410] + MEM[38451];
assign MEM[44137] = MEM[38412] + MEM[38487];
assign MEM[44138] = MEM[38417] + MEM[38471];
assign MEM[44139] = MEM[38421] + MEM[38464];
assign MEM[44140] = MEM[38422] + MEM[38480];
assign MEM[44141] = MEM[38424] + MEM[38458];
assign MEM[44142] = MEM[38425] + MEM[38460];
assign MEM[44143] = MEM[38428] + MEM[38496];
assign MEM[44144] = MEM[38430] + MEM[38504];
assign MEM[44145] = MEM[38432] + MEM[38508];
assign MEM[44146] = MEM[38433] + MEM[38549];
assign MEM[44147] = MEM[38434] + MEM[38494];
assign MEM[44148] = MEM[38436] + MEM[38529];
assign MEM[44149] = MEM[38437] + MEM[38501];
assign MEM[44150] = MEM[38438] + MEM[38474];
assign MEM[44151] = MEM[38439] + MEM[38482];
assign MEM[44152] = MEM[38440] + MEM[38531];
assign MEM[44153] = MEM[38441] + MEM[38462];
assign MEM[44154] = MEM[38442] + MEM[38489];
assign MEM[44155] = MEM[38444] + MEM[38466];
assign MEM[44156] = MEM[38445] + MEM[38486];
assign MEM[44157] = MEM[38447] + MEM[38470];
assign MEM[44158] = MEM[38449] + MEM[38461];
assign MEM[44159] = MEM[38450] + MEM[38593];
assign MEM[44160] = MEM[38453] + MEM[38560];
assign MEM[44161] = MEM[38454] + MEM[38497];
assign MEM[44162] = MEM[38455] + MEM[38520];
assign MEM[44163] = MEM[38456] + MEM[38476];
assign MEM[44164] = MEM[38459] + MEM[38523];
assign MEM[44165] = MEM[38463] + MEM[38495];
assign MEM[44166] = MEM[38465] + MEM[38557];
assign MEM[44167] = MEM[38469] + MEM[38574];
assign MEM[44168] = MEM[38472] + MEM[38533];
assign MEM[44169] = MEM[38475] + MEM[38589];
assign MEM[44170] = MEM[38477] + MEM[38658];
assign MEM[44171] = MEM[38478] + MEM[38493];
assign MEM[44172] = MEM[38479] + MEM[38567];
assign MEM[44173] = MEM[38481] + MEM[38583];
assign MEM[44174] = MEM[38484] + MEM[38555];
assign MEM[44175] = MEM[38485] + MEM[38548];
assign MEM[44176] = MEM[38488] + MEM[38566];
assign MEM[44177] = MEM[38490] + MEM[38610];
assign MEM[44178] = MEM[38491] + MEM[38521];
assign MEM[44179] = MEM[38492] + MEM[38516];
assign MEM[44180] = MEM[38499] + MEM[38685];
assign MEM[44181] = MEM[38500] + MEM[38617];
assign MEM[44182] = MEM[38502] + MEM[38608];
assign MEM[44183] = MEM[38503] + MEM[38539];
assign MEM[44184] = MEM[38505] + MEM[38538];
assign MEM[44185] = MEM[38506] + MEM[38661];
assign MEM[44186] = MEM[38507] + MEM[38542];
assign MEM[44187] = MEM[38509] + MEM[38629];
assign MEM[44188] = MEM[38510] + MEM[38632];
assign MEM[44189] = MEM[38511] + MEM[38599];
assign MEM[44190] = MEM[38512] + MEM[38598];
assign MEM[44191] = MEM[38513] + MEM[38570];
assign MEM[44192] = MEM[38514] + MEM[38619];
assign MEM[44193] = MEM[38515] + MEM[38534];
assign MEM[44194] = MEM[38518] + MEM[38535];
assign MEM[44195] = MEM[38519] + MEM[38587];
assign MEM[44196] = MEM[38524] + MEM[38550];
assign MEM[44197] = MEM[38525] + MEM[38719];
assign MEM[44198] = MEM[38526] + MEM[38573];
assign MEM[44199] = MEM[38527] + MEM[38591];
assign MEM[44200] = MEM[38528] + MEM[38607];
assign MEM[44201] = MEM[38530] + MEM[38578];
assign MEM[44202] = MEM[38532] + MEM[38551];
assign MEM[44203] = MEM[38536] + MEM[38558];
assign MEM[44204] = MEM[38537] + MEM[38577];
assign MEM[44205] = MEM[38540] + MEM[38563];
assign MEM[44206] = MEM[38541] + MEM[38623];
assign MEM[44207] = MEM[38544] + MEM[38595];
assign MEM[44208] = MEM[38545] + MEM[38559];
assign MEM[44209] = MEM[38546] + MEM[38672];
assign MEM[44210] = MEM[38547] + MEM[38588];
assign MEM[44211] = MEM[38552] + MEM[38576];
assign MEM[44212] = MEM[38553] + MEM[38568];
assign MEM[44213] = MEM[38554] + MEM[38611];
assign MEM[44214] = MEM[38556] + MEM[38652];
assign MEM[44215] = MEM[38561] + MEM[38592];
assign MEM[44216] = MEM[38562] + MEM[38637];
assign MEM[44217] = MEM[38564] + MEM[38596];
assign MEM[44218] = MEM[38565] + MEM[38668];
assign MEM[44219] = MEM[38569] + MEM[38605];
assign MEM[44220] = MEM[38571] + MEM[38670];
assign MEM[44221] = MEM[38572] + MEM[38600];
assign MEM[44222] = MEM[38575] + MEM[38620];
assign MEM[44223] = MEM[38579] + MEM[38634];
assign MEM[44224] = MEM[38580] + MEM[38676];
assign MEM[44225] = MEM[38581] + MEM[38602];
assign MEM[44226] = MEM[38582] + MEM[38631];
assign MEM[44227] = MEM[38584] + MEM[38678];
assign MEM[44228] = MEM[38585] + MEM[38681];
assign MEM[44229] = MEM[38586] + MEM[38606];
assign MEM[44230] = MEM[38590] + MEM[38613];
assign MEM[44231] = MEM[38594] + MEM[38642];
assign MEM[44232] = MEM[38597] + MEM[38666];
assign MEM[44233] = MEM[38601] + MEM[38643];
assign MEM[44234] = MEM[38603] + MEM[38707];
assign MEM[44235] = MEM[38604] + MEM[38674];
assign MEM[44236] = MEM[38609] + MEM[38625];
assign MEM[44237] = MEM[38612] + MEM[38679];
assign MEM[44238] = MEM[38614] + MEM[38677];
assign MEM[44239] = MEM[38615] + MEM[38635];
assign MEM[44240] = MEM[38616] + MEM[38651];
assign MEM[44241] = MEM[38618] + MEM[38694];
assign MEM[44242] = MEM[38621] + MEM[38682];
assign MEM[44243] = MEM[38622] + MEM[38671];
assign MEM[44244] = MEM[38624] + MEM[38698];
assign MEM[44245] = MEM[38626] + MEM[38646];
assign MEM[44246] = MEM[38627] + MEM[38691];
assign MEM[44247] = MEM[38628] + MEM[38683];
assign MEM[44248] = MEM[38630] + MEM[38709];
assign MEM[44249] = MEM[38633] + MEM[38695];
assign MEM[44250] = MEM[38636] + MEM[38704];
assign MEM[44251] = MEM[38638] + MEM[38703];
assign MEM[44252] = MEM[38639] + MEM[38706];
assign MEM[44253] = MEM[38640] + MEM[38715];
assign MEM[44254] = MEM[38641] + MEM[38696];
assign MEM[44255] = MEM[38644] + MEM[38657];
assign MEM[44256] = MEM[38645] + MEM[38767];
assign MEM[44257] = MEM[38647] + MEM[38687];
assign MEM[44258] = MEM[38648] + MEM[38675];
assign MEM[44259] = MEM[38649] + MEM[38733];
assign MEM[44260] = MEM[38650] + MEM[38690];
assign MEM[44261] = MEM[38653] + MEM[38686];
assign MEM[44262] = MEM[38654] + MEM[38772];
assign MEM[44263] = MEM[38655] + MEM[38769];
assign MEM[44264] = MEM[38656] + MEM[38913];
assign MEM[44265] = MEM[38659] + MEM[38701];
assign MEM[44266] = MEM[38660] + MEM[38725];
assign MEM[44267] = MEM[38662] + MEM[38788];
assign MEM[44268] = MEM[38663] + MEM[38689];
assign MEM[44269] = MEM[38664] + MEM[38740];
assign MEM[44270] = MEM[38665] + MEM[38705];
assign MEM[44271] = MEM[38667] + MEM[38768];
assign MEM[44272] = MEM[38669] + MEM[38766];
assign MEM[44273] = MEM[38673] + MEM[38799];
assign MEM[44274] = MEM[38680] + MEM[38724];
assign MEM[44275] = MEM[38684] + MEM[38801];
assign MEM[44276] = MEM[38688] + MEM[38729];
assign MEM[44277] = MEM[38692] + MEM[38714];
assign MEM[44278] = MEM[38693] + MEM[38712];
assign MEM[44279] = MEM[38697] + MEM[38782];
assign MEM[44280] = MEM[38699] + MEM[38722];
assign MEM[44281] = MEM[38700] + MEM[38762];
assign MEM[44282] = MEM[38702] + MEM[38770];
assign MEM[44283] = MEM[38708] + MEM[38850];
assign MEM[44284] = MEM[38710] + MEM[38739];
assign MEM[44285] = MEM[38711] + MEM[38745];
assign MEM[44286] = MEM[38713] + MEM[38804];
assign MEM[44287] = MEM[38716] + MEM[38747];
assign MEM[44288] = MEM[38717] + MEM[38781];
assign MEM[44289] = MEM[38718] + MEM[38752];
assign MEM[44290] = MEM[38720] + MEM[38761];
assign MEM[44291] = MEM[38721] + MEM[38754];
assign MEM[44292] = MEM[38723] + MEM[38855];
assign MEM[44293] = MEM[38726] + MEM[38771];
assign MEM[44294] = MEM[38727] + MEM[38778];
assign MEM[44295] = MEM[38728] + MEM[38811];
assign MEM[44296] = MEM[38730] + MEM[38744];
assign MEM[44297] = MEM[38731] + MEM[38883];
assign MEM[44298] = MEM[38732] + MEM[38755];
assign MEM[44299] = MEM[38734] + MEM[38821];
assign MEM[44300] = MEM[38735] + MEM[38742];
assign MEM[44301] = MEM[38736] + MEM[38806];
assign MEM[44302] = MEM[38737] + MEM[38774];
assign MEM[44303] = MEM[38738] + MEM[38870];
assign MEM[44304] = MEM[38741] + MEM[38810];
assign MEM[44305] = MEM[38743] + MEM[38758];
assign MEM[44306] = MEM[38746] + MEM[38924];
assign MEM[44307] = MEM[38748] + MEM[38798];
assign MEM[44308] = MEM[38749] + MEM[38780];
assign MEM[44309] = MEM[38750] + MEM[38818];
assign MEM[44310] = MEM[38751] + MEM[38854];
assign MEM[44311] = MEM[38753] + MEM[38819];
assign MEM[44312] = MEM[38756] + MEM[38807];
assign MEM[44313] = MEM[38757] + MEM[38792];
assign MEM[44314] = MEM[38759] + MEM[38824];
assign MEM[44315] = MEM[38760] + MEM[38859];
assign MEM[44316] = MEM[38763] + MEM[38872];
assign MEM[44317] = MEM[38764] + MEM[38779];
assign MEM[44318] = MEM[38765] + MEM[38783];
assign MEM[44319] = MEM[38773] + MEM[38828];
assign MEM[44320] = MEM[38775] + MEM[38790];
assign MEM[44321] = MEM[38776] + MEM[38833];
assign MEM[44322] = MEM[38777] + MEM[38791];
assign MEM[44323] = MEM[38784] + MEM[38939];
assign MEM[44324] = MEM[38785] + MEM[38823];
assign MEM[44325] = MEM[38786] + MEM[38812];
assign MEM[44326] = MEM[38787] + MEM[38955];
assign MEM[44327] = MEM[38789] + MEM[38803];
assign MEM[44328] = MEM[38793] + MEM[38829];
assign MEM[44329] = MEM[38794] + MEM[38864];
assign MEM[44330] = MEM[38795] + MEM[38839];
assign MEM[44331] = MEM[38796] + MEM[38834];
assign MEM[44332] = MEM[38797] + MEM[38931];
assign MEM[44333] = MEM[38800] + MEM[38861];
assign MEM[44334] = MEM[38802] + MEM[38835];
assign MEM[44335] = MEM[38805] + MEM[38830];
assign MEM[44336] = MEM[38808] + MEM[38841];
assign MEM[44337] = MEM[38809] + MEM[38820];
assign MEM[44338] = MEM[38813] + MEM[38837];
assign MEM[44339] = MEM[38814] + MEM[38826];
assign MEM[44340] = MEM[38815] + MEM[38866];
assign MEM[44341] = MEM[38816] + MEM[38863];
assign MEM[44342] = MEM[38817] + MEM[38845];
assign MEM[44343] = MEM[38822] + MEM[38896];
assign MEM[44344] = MEM[38825] + MEM[38880];
assign MEM[44345] = MEM[38827] + MEM[38851];
assign MEM[44346] = MEM[38831] + MEM[38949];
assign MEM[44347] = MEM[38832] + MEM[39045];
assign MEM[44348] = MEM[38836] + MEM[38969];
assign MEM[44349] = MEM[38838] + MEM[38874];
assign MEM[44350] = MEM[38840] + MEM[38871];
assign MEM[44351] = MEM[38842] + MEM[38858];
assign MEM[44352] = MEM[38843] + MEM[38865];
assign MEM[44353] = MEM[38844] + MEM[38954];
assign MEM[44354] = MEM[38846] + MEM[38882];
assign MEM[44355] = MEM[38847] + MEM[38884];
assign MEM[44356] = MEM[38848] + MEM[38894];
assign MEM[44357] = MEM[38849] + MEM[38878];
assign MEM[44358] = MEM[38852] + MEM[38886];
assign MEM[44359] = MEM[38853] + MEM[38901];
assign MEM[44360] = MEM[38856] + MEM[38947];
assign MEM[44361] = MEM[38857] + MEM[38899];
assign MEM[44362] = MEM[38860] + MEM[38933];
assign MEM[44363] = MEM[38862] + MEM[38885];
assign MEM[44364] = MEM[38867] + MEM[38891];
assign MEM[44365] = MEM[38868] + MEM[39090];
assign MEM[44366] = MEM[38869] + MEM[38915];
assign MEM[44367] = MEM[38873] + MEM[38950];
assign MEM[44368] = MEM[38875] + MEM[38905];
assign MEM[44369] = MEM[38876] + MEM[38957];
assign MEM[44370] = MEM[38877] + MEM[38916];
assign MEM[44371] = MEM[38879] + MEM[38895];
assign MEM[44372] = MEM[38881] + MEM[38923];
assign MEM[44373] = MEM[38887] + MEM[38928];
assign MEM[44374] = MEM[38888] + MEM[38900];
assign MEM[44375] = MEM[38889] + MEM[38946];
assign MEM[44376] = MEM[38890] + MEM[38945];
assign MEM[44377] = MEM[38892] + MEM[38951];
assign MEM[44378] = MEM[38893] + MEM[38962];
assign MEM[44379] = MEM[38897] + MEM[38919];
assign MEM[44380] = MEM[38898] + MEM[38912];
assign MEM[44381] = MEM[38902] + MEM[38991];
assign MEM[44382] = MEM[38903] + MEM[38922];
assign MEM[44383] = MEM[38904] + MEM[38956];
assign MEM[44384] = MEM[38906] + MEM[39085];
assign MEM[44385] = MEM[38907] + MEM[38970];
assign MEM[44386] = MEM[38908] + MEM[38964];
assign MEM[44387] = MEM[38909] + MEM[38942];
assign MEM[44388] = MEM[38910] + MEM[38925];
assign MEM[44389] = MEM[38911] + MEM[38998];
assign MEM[44390] = MEM[38914] + MEM[38963];
assign MEM[44391] = MEM[38917] + MEM[38952];
assign MEM[44392] = MEM[38918] + MEM[39028];
assign MEM[44393] = MEM[38920] + MEM[38959];
assign MEM[44394] = MEM[38921] + MEM[39065];
assign MEM[44395] = MEM[38926] + MEM[38993];
assign MEM[44396] = MEM[38927] + MEM[38938];
assign MEM[44397] = MEM[38929] + MEM[38987];
assign MEM[44398] = MEM[38930] + MEM[38976];
assign MEM[44399] = MEM[38932] + MEM[38977];
assign MEM[44400] = MEM[38934] + MEM[38967];
assign MEM[44401] = MEM[38935] + MEM[39005];
assign MEM[44402] = MEM[38936] + MEM[38973];
assign MEM[44403] = MEM[38937] + MEM[39008];
assign MEM[44404] = MEM[38940] + MEM[39012];
assign MEM[44405] = MEM[38941] + MEM[39040];
assign MEM[44406] = MEM[38943] + MEM[39018];
assign MEM[44407] = MEM[38944] + MEM[39039];
assign MEM[44408] = MEM[38948] + MEM[39000];
assign MEM[44409] = MEM[38953] + MEM[39027];
assign MEM[44410] = MEM[38958] + MEM[39002];
assign MEM[44411] = MEM[38960] + MEM[38986];
assign MEM[44412] = MEM[38961] + MEM[39006];
assign MEM[44413] = MEM[38965] + MEM[39062];
assign MEM[44414] = MEM[38966] + MEM[39060];
assign MEM[44415] = MEM[38968] + MEM[39029];
assign MEM[44416] = MEM[38971] + MEM[38997];
assign MEM[44417] = MEM[38972] + MEM[39001];
assign MEM[44418] = MEM[38974] + MEM[39020];
assign MEM[44419] = MEM[38975] + MEM[38989];
assign MEM[44420] = MEM[38978] + MEM[39013];
assign MEM[44421] = MEM[38979] + MEM[39016];
assign MEM[44422] = MEM[38980] + MEM[39017];
assign MEM[44423] = MEM[38981] + MEM[39056];
assign MEM[44424] = MEM[38982] + MEM[39023];
assign MEM[44425] = MEM[38983] + MEM[39089];
assign MEM[44426] = MEM[38984] + MEM[39066];
assign MEM[44427] = MEM[38985] + MEM[39136];
assign MEM[44428] = MEM[38988] + MEM[39084];
assign MEM[44429] = MEM[38990] + MEM[39003];
assign MEM[44430] = MEM[38992] + MEM[39098];
assign MEM[44431] = MEM[38994] + MEM[39081];
assign MEM[44432] = MEM[38995] + MEM[39058];
assign MEM[44433] = MEM[38996] + MEM[39113];
assign MEM[44434] = MEM[38999] + MEM[39021];
assign MEM[44435] = MEM[39004] + MEM[39051];
assign MEM[44436] = MEM[39007] + MEM[39091];
assign MEM[44437] = MEM[39009] + MEM[39139];
assign MEM[44438] = MEM[39010] + MEM[39049];
assign MEM[44439] = MEM[39011] + MEM[39116];
assign MEM[44440] = MEM[39014] + MEM[39052];
assign MEM[44441] = MEM[39015] + MEM[39188];
assign MEM[44442] = MEM[39019] + MEM[39044];
assign MEM[44443] = MEM[39022] + MEM[39104];
assign MEM[44444] = MEM[39024] + MEM[39041];
assign MEM[44445] = MEM[39025] + MEM[39122];
assign MEM[44446] = MEM[39026] + MEM[39037];
assign MEM[44447] = MEM[39030] + MEM[39043];
assign MEM[44448] = MEM[39031] + MEM[39102];
assign MEM[44449] = MEM[39032] + MEM[39174];
assign MEM[44450] = MEM[39033] + MEM[39095];
assign MEM[44451] = MEM[39034] + MEM[39201];
assign MEM[44452] = MEM[39035] + MEM[39169];
assign MEM[44453] = MEM[39036] + MEM[39141];
assign MEM[44454] = MEM[39038] + MEM[39072];
assign MEM[44455] = MEM[39042] + MEM[39115];
assign MEM[44456] = MEM[39046] + MEM[39107];
assign MEM[44457] = MEM[39047] + MEM[39118];
assign MEM[44458] = MEM[39048] + MEM[39082];
assign MEM[44459] = MEM[39050] + MEM[39092];
assign MEM[44460] = MEM[39053] + MEM[39055];
assign MEM[44461] = MEM[39054] + MEM[39167];
assign MEM[44462] = MEM[39057] + MEM[39105];
assign MEM[44463] = MEM[39059] + MEM[39078];
assign MEM[44464] = MEM[39061] + MEM[39150];
assign MEM[44465] = MEM[39063] + MEM[39087];
assign MEM[44466] = MEM[39064] + MEM[39209];
assign MEM[44467] = MEM[39067] + MEM[39147];
assign MEM[44468] = MEM[39068] + MEM[39153];
assign MEM[44469] = MEM[39069] + MEM[39121];
assign MEM[44470] = MEM[39070] + MEM[39114];
assign MEM[44471] = MEM[39071] + MEM[39086];
assign MEM[44472] = MEM[39073] + MEM[39160];
assign MEM[44473] = MEM[39074] + MEM[39158];
assign MEM[44474] = MEM[39075] + MEM[39163];
assign MEM[44475] = MEM[39076] + MEM[39119];
assign MEM[44476] = MEM[39077] + MEM[39146];
assign MEM[44477] = MEM[39079] + MEM[39125];
assign MEM[44478] = MEM[39080] + MEM[39096];
assign MEM[44479] = MEM[39083] + MEM[39142];
assign MEM[44480] = MEM[39088] + MEM[39140];
assign MEM[44481] = MEM[39093] + MEM[39109];
assign MEM[44482] = MEM[39094] + MEM[39355];
assign MEM[44483] = MEM[39097] + MEM[39144];
assign MEM[44484] = MEM[39099] + MEM[39128];
assign MEM[44485] = MEM[39100] + MEM[39149];
assign MEM[44486] = MEM[39101] + MEM[39195];
assign MEM[44487] = MEM[39103] + MEM[39213];
assign MEM[44488] = MEM[39106] + MEM[39198];
assign MEM[44489] = MEM[39108] + MEM[39145];
assign MEM[44490] = MEM[39110] + MEM[39129];
assign MEM[44491] = MEM[39111] + MEM[39159];
assign MEM[44492] = MEM[39112] + MEM[39176];
assign MEM[44493] = MEM[39117] + MEM[39148];
assign MEM[44494] = MEM[39120] + MEM[39184];
assign MEM[44495] = MEM[39123] + MEM[39164];
assign MEM[44496] = MEM[39124] + MEM[39132];
assign MEM[44497] = MEM[39126] + MEM[39200];
assign MEM[44498] = MEM[39127] + MEM[39227];
assign MEM[44499] = MEM[39130] + MEM[39170];
assign MEM[44500] = MEM[39131] + MEM[39199];
assign MEM[44501] = MEM[39133] + MEM[39313];
assign MEM[44502] = MEM[39134] + MEM[39154];
assign MEM[44503] = MEM[39135] + MEM[39168];
assign MEM[44504] = MEM[39137] + MEM[39151];
assign MEM[44505] = MEM[39138] + MEM[39191];
assign MEM[44506] = MEM[39143] + MEM[39289];
assign MEM[44507] = MEM[39152] + MEM[39306];
assign MEM[44508] = MEM[39155] + MEM[39202];
assign MEM[44509] = MEM[39156] + MEM[39192];
assign MEM[44510] = MEM[39157] + MEM[39248];
assign MEM[44511] = MEM[39161] + MEM[39312];
assign MEM[44512] = MEM[39162] + MEM[39182];
assign MEM[44513] = MEM[39165] + MEM[39242];
assign MEM[44514] = MEM[39166] + MEM[39240];
assign MEM[44515] = MEM[39171] + MEM[39215];
assign MEM[44516] = MEM[39172] + MEM[39212];
assign MEM[44517] = MEM[39173] + MEM[39224];
assign MEM[44518] = MEM[39175] + MEM[39262];
assign MEM[44519] = MEM[39177] + MEM[39222];
assign MEM[44520] = MEM[39178] + MEM[39230];
assign MEM[44521] = MEM[39179] + MEM[39204];
assign MEM[44522] = MEM[39180] + MEM[39279];
assign MEM[44523] = MEM[39181] + MEM[39270];
assign MEM[44524] = MEM[39183] + MEM[39203];
assign MEM[44525] = MEM[39185] + MEM[39214];
assign MEM[44526] = MEM[39186] + MEM[39318];
assign MEM[44527] = MEM[39187] + MEM[39239];
assign MEM[44528] = MEM[39189] + MEM[39283];
assign MEM[44529] = MEM[39190] + MEM[39228];
assign MEM[44530] = MEM[39193] + MEM[39345];
assign MEM[44531] = MEM[39194] + MEM[39253];
assign MEM[44532] = MEM[39196] + MEM[39237];
assign MEM[44533] = MEM[39197] + MEM[39267];
assign MEM[44534] = MEM[39205] + MEM[39216];
assign MEM[44535] = MEM[39206] + MEM[39298];
assign MEM[44536] = MEM[39207] + MEM[39285];
assign MEM[44537] = MEM[39208] + MEM[39243];
assign MEM[44538] = MEM[39210] + MEM[39309];
assign MEM[44539] = MEM[39211] + MEM[39235];
assign MEM[44540] = MEM[39217] + MEM[39256];
assign MEM[44541] = MEM[39218] + MEM[39315];
assign MEM[44542] = MEM[39219] + MEM[39303];
assign MEM[44543] = MEM[39220] + MEM[39308];
assign MEM[44544] = MEM[39221] + MEM[39260];
assign MEM[44545] = MEM[39223] + MEM[39244];
assign MEM[44546] = MEM[39225] + MEM[39422];
assign MEM[44547] = MEM[39226] + MEM[39282];
assign MEM[44548] = MEM[39229] + MEM[39442];
assign MEM[44549] = MEM[39231] + MEM[39343];
assign MEM[44550] = MEM[39232] + MEM[39261];
assign MEM[44551] = MEM[39233] + MEM[39372];
assign MEM[44552] = MEM[39234] + MEM[39292];
assign MEM[44553] = MEM[39236] + MEM[39326];
assign MEM[44554] = MEM[39238] + MEM[39288];
assign MEM[44555] = MEM[39241] + MEM[39264];
assign MEM[44556] = MEM[39245] + MEM[39259];
assign MEM[44557] = MEM[39246] + MEM[39296];
assign MEM[44558] = MEM[39247] + MEM[39344];
assign MEM[44559] = MEM[39249] + MEM[39378];
assign MEM[44560] = MEM[39250] + MEM[39356];
assign MEM[44561] = MEM[39251] + MEM[39278];
assign MEM[44562] = MEM[39252] + MEM[39330];
assign MEM[44563] = MEM[39254] + MEM[39363];
assign MEM[44564] = MEM[39255] + MEM[39277];
assign MEM[44565] = MEM[39257] + MEM[39302];
assign MEM[44566] = MEM[39258] + MEM[39393];
assign MEM[44567] = MEM[39263] + MEM[39294];
assign MEM[44568] = MEM[39265] + MEM[39336];
assign MEM[44569] = MEM[39266] + MEM[39291];
assign MEM[44570] = MEM[39268] + MEM[39319];
assign MEM[44571] = MEM[39269] + MEM[39320];
assign MEM[44572] = MEM[39271] + MEM[39293];
assign MEM[44573] = MEM[39272] + MEM[39299];
assign MEM[44574] = MEM[39273] + MEM[39370];
assign MEM[44575] = MEM[39274] + MEM[39390];
assign MEM[44576] = MEM[39275] + MEM[39280];
assign MEM[44577] = MEM[39276] + MEM[39383];
assign MEM[44578] = MEM[39281] + MEM[39365];
assign MEM[44579] = MEM[39284] + MEM[39301];
assign MEM[44580] = MEM[39286] + MEM[39413];
assign MEM[44581] = MEM[39287] + MEM[39399];
assign MEM[44582] = MEM[39290] + MEM[39337];
assign MEM[44583] = MEM[39295] + MEM[39340];
assign MEM[44584] = MEM[39297] + MEM[39436];
assign MEM[44585] = MEM[39300] + MEM[39428];
assign MEM[44586] = MEM[39304] + MEM[39368];
assign MEM[44587] = MEM[39305] + MEM[39317];
assign MEM[44588] = MEM[39307] + MEM[39325];
assign MEM[44589] = MEM[39310] + MEM[39341];
assign MEM[44590] = MEM[39311] + MEM[39351];
assign MEM[44591] = MEM[39314] + MEM[39354];
assign MEM[44592] = MEM[39316] + MEM[39366];
assign MEM[44593] = MEM[39321] + MEM[39342];
assign MEM[44594] = MEM[39322] + MEM[39402];
assign MEM[44595] = MEM[39323] + MEM[39361];
assign MEM[44596] = MEM[39324] + MEM[39380];
assign MEM[44597] = MEM[39327] + MEM[39525];
assign MEM[44598] = MEM[39328] + MEM[39353];
assign MEM[44599] = MEM[39329] + MEM[39421];
assign MEM[44600] = MEM[39331] + MEM[39431];
assign MEM[44601] = MEM[39332] + MEM[39387];
assign MEM[44602] = MEM[39333] + MEM[39369];
assign MEM[44603] = MEM[39334] + MEM[39448];
assign MEM[44604] = MEM[39335] + MEM[39417];
assign MEM[44605] = MEM[39338] + MEM[39359];
assign MEM[44606] = MEM[39339] + MEM[39374];
assign MEM[44607] = MEM[39346] + MEM[39411];
assign MEM[44608] = MEM[39347] + MEM[39501];
assign MEM[44609] = MEM[39348] + MEM[39521];
assign MEM[44610] = MEM[39349] + MEM[39388];
assign MEM[44611] = MEM[39350] + MEM[39391];
assign MEM[44612] = MEM[39352] + MEM[39382];
assign MEM[44613] = MEM[39357] + MEM[39561];
assign MEM[44614] = MEM[39358] + MEM[39415];
assign MEM[44615] = MEM[39360] + MEM[39416];
assign MEM[44616] = MEM[39362] + MEM[39454];
assign MEM[44617] = MEM[39364] + MEM[39494];
assign MEM[44618] = MEM[39367] + MEM[39445];
assign MEM[44619] = MEM[39371] + MEM[39401];
assign MEM[44620] = MEM[39373] + MEM[39435];
assign MEM[44621] = MEM[39375] + MEM[39377];
assign MEM[44622] = MEM[39376] + MEM[39394];
assign MEM[44623] = MEM[39379] + MEM[39423];
assign MEM[44624] = MEM[39381] + MEM[39427];
assign MEM[44625] = MEM[39384] + MEM[39464];
assign MEM[44626] = MEM[39385] + MEM[39472];
assign MEM[44627] = MEM[39386] + MEM[39434];
assign MEM[44628] = MEM[39389] + MEM[39404];
assign MEM[44629] = MEM[39392] + MEM[39455];
assign MEM[44630] = MEM[39395] + MEM[39470];
assign MEM[44631] = MEM[39396] + MEM[39429];
assign MEM[44632] = MEM[39397] + MEM[39426];
assign MEM[44633] = MEM[39398] + MEM[39412];
assign MEM[44634] = MEM[39400] + MEM[39410];
assign MEM[44635] = MEM[39403] + MEM[39513];
assign MEM[44636] = MEM[39405] + MEM[39511];
assign MEM[44637] = MEM[39406] + MEM[39439];
assign MEM[44638] = MEM[39407] + MEM[39465];
assign MEM[44639] = MEM[39408] + MEM[39419];
assign MEM[44640] = MEM[39409] + MEM[39507];
assign MEM[44641] = MEM[39414] + MEM[39460];
assign MEM[44642] = MEM[39418] + MEM[39481];
assign MEM[44643] = MEM[39420] + MEM[39450];
assign MEM[44644] = MEM[39424] + MEM[39512];
assign MEM[44645] = MEM[39425] + MEM[39473];
assign MEM[44646] = MEM[39430] + MEM[39443];
assign MEM[44647] = MEM[39432] + MEM[39468];
assign MEM[44648] = MEM[39433] + MEM[39447];
assign MEM[44649] = MEM[39437] + MEM[39471];
assign MEM[44650] = MEM[39438] + MEM[39484];
assign MEM[44651] = MEM[39440] + MEM[39497];
assign MEM[44652] = MEM[39441] + MEM[39563];
assign MEM[44653] = MEM[39444] + MEM[39491];
assign MEM[44654] = MEM[39446] + MEM[39503];
assign MEM[44655] = MEM[39449] + MEM[39546];
assign MEM[44656] = MEM[39451] + MEM[39489];
assign MEM[44657] = MEM[39452] + MEM[39492];
assign MEM[44658] = MEM[39453] + MEM[39540];
assign MEM[44659] = MEM[39456] + MEM[39573];
assign MEM[44660] = MEM[39457] + MEM[39534];
assign MEM[44661] = MEM[39458] + MEM[39495];
assign MEM[44662] = MEM[39459] + MEM[39524];
assign MEM[44663] = MEM[39461] + MEM[39477];
assign MEM[44664] = MEM[39462] + MEM[39500];
assign MEM[44665] = MEM[39463] + MEM[39516];
assign MEM[44666] = MEM[39466] + MEM[39564];
assign MEM[44667] = MEM[39467] + MEM[39508];
assign MEM[44668] = MEM[39469] + MEM[39493];
assign MEM[44669] = MEM[39474] + MEM[39483];
assign MEM[44670] = MEM[39475] + MEM[39515];
assign MEM[44671] = MEM[39476] + MEM[39633];
assign MEM[44672] = MEM[39478] + MEM[39502];
assign MEM[44673] = MEM[39479] + MEM[39642];
assign MEM[44674] = MEM[39480] + MEM[39490];
assign MEM[44675] = MEM[39482] + MEM[39499];
assign MEM[44676] = MEM[39485] + MEM[39555];
assign MEM[44677] = MEM[39486] + MEM[39577];
assign MEM[44678] = MEM[39487] + MEM[39599];
assign MEM[44679] = MEM[39488] + MEM[39571];
assign MEM[44680] = MEM[39496] + MEM[39541];
assign MEM[44681] = MEM[39498] + MEM[39532];
assign MEM[44682] = MEM[39504] + MEM[39613];
assign MEM[44683] = MEM[39505] + MEM[39539];
assign MEM[44684] = MEM[39506] + MEM[39543];
assign MEM[44685] = MEM[39509] + MEM[39568];
assign MEM[44686] = MEM[39510] + MEM[39560];
assign MEM[44687] = MEM[39514] + MEM[39569];
assign MEM[44688] = MEM[39517] + MEM[39616];
assign MEM[44689] = MEM[39518] + MEM[39547];
assign MEM[44690] = MEM[39519] + MEM[39558];
assign MEM[44691] = MEM[39520] + MEM[39621];
assign MEM[44692] = MEM[39522] + MEM[39550];
assign MEM[44693] = MEM[39523] + MEM[39582];
assign MEM[44694] = MEM[39526] + MEM[39585];
assign MEM[44695] = MEM[39527] + MEM[39590];
assign MEM[44696] = MEM[39528] + MEM[39622];
assign MEM[44697] = MEM[39529] + MEM[39570];
assign MEM[44698] = MEM[39530] + MEM[39612];
assign MEM[44699] = MEM[39531] + MEM[39565];
assign MEM[44700] = MEM[39533] + MEM[39614];
assign MEM[44701] = MEM[39535] + MEM[39580];
assign MEM[44702] = MEM[39536] + MEM[39594];
assign MEM[44703] = MEM[39537] + MEM[39566];
assign MEM[44704] = MEM[39538] + MEM[39592];
assign MEM[44705] = MEM[39542] + MEM[39587];
assign MEM[44706] = MEM[39544] + MEM[39617];
assign MEM[44707] = MEM[39545] + MEM[39615];
assign MEM[44708] = MEM[39548] + MEM[39576];
assign MEM[44709] = MEM[39549] + MEM[39624];
assign MEM[44710] = MEM[39551] + MEM[39749];
assign MEM[44711] = MEM[39552] + MEM[39602];
assign MEM[44712] = MEM[39553] + MEM[39601];
assign MEM[44713] = MEM[39554] + MEM[39625];
assign MEM[44714] = MEM[39556] + MEM[39655];
assign MEM[44715] = MEM[39557] + MEM[39727];
assign MEM[44716] = MEM[39559] + MEM[39668];
assign MEM[44717] = MEM[39562] + MEM[39595];
assign MEM[44718] = MEM[39567] + MEM[39628];
assign MEM[44719] = MEM[39572] + MEM[39654];
assign MEM[44720] = MEM[39574] + MEM[39631];
assign MEM[44721] = MEM[39575] + MEM[39726];
assign MEM[44722] = MEM[39578] + MEM[39623];
assign MEM[44723] = MEM[39579] + MEM[39672];
assign MEM[44724] = MEM[39581] + MEM[39603];
assign MEM[44725] = MEM[39583] + MEM[39667];
assign MEM[44726] = MEM[39584] + MEM[39604];
assign MEM[44727] = MEM[39586] + MEM[39678];
assign MEM[44728] = MEM[39588] + MEM[39653];
assign MEM[44729] = MEM[39589] + MEM[39619];
assign MEM[44730] = MEM[39591] + MEM[39673];
assign MEM[44731] = MEM[39593] + MEM[39659];
assign MEM[44732] = MEM[39596] + MEM[39664];
assign MEM[44733] = MEM[39597] + MEM[39632];
assign MEM[44734] = MEM[39598] + MEM[39644];
assign MEM[44735] = MEM[39600] + MEM[39641];
assign MEM[44736] = MEM[39605] + MEM[39650];
assign MEM[44737] = MEM[39606] + MEM[39647];
assign MEM[44738] = MEM[39607] + MEM[39652];
assign MEM[44739] = MEM[39608] + MEM[39638];
assign MEM[44740] = MEM[39609] + MEM[39677];
assign MEM[44741] = MEM[39610] + MEM[39688];
assign MEM[44742] = MEM[39611] + MEM[39696];
assign MEM[44743] = MEM[39618] + MEM[39656];
assign MEM[44744] = MEM[39620] + MEM[39637];
assign MEM[44745] = MEM[39626] + MEM[39720];
assign MEM[44746] = MEM[39627] + MEM[39643];
assign MEM[44747] = MEM[39629] + MEM[39689];
assign MEM[44748] = MEM[39630] + MEM[39759];
assign MEM[44749] = MEM[39634] + MEM[39636];
assign MEM[44750] = MEM[39635] + MEM[39836];
assign MEM[44751] = MEM[39639] + MEM[39695];
assign MEM[44752] = MEM[39640] + MEM[39674];
assign MEM[44753] = MEM[39645] + MEM[39666];
assign MEM[44754] = MEM[39646] + MEM[39706];
assign MEM[44755] = MEM[39648] + MEM[39703];
assign MEM[44756] = MEM[39649] + MEM[39795];
assign MEM[44757] = MEM[39651] + MEM[39661];
assign MEM[44758] = MEM[39657] + MEM[39710];
assign MEM[44759] = MEM[39658] + MEM[39760];
assign MEM[44760] = MEM[39660] + MEM[39690];
assign MEM[44761] = MEM[39662] + MEM[39685];
assign MEM[44762] = MEM[39663] + MEM[39698];
assign MEM[44763] = MEM[39665] + MEM[39715];
assign MEM[44764] = MEM[39669] + MEM[39693];
assign MEM[44765] = MEM[39670] + MEM[39716];
assign MEM[44766] = MEM[39671] + MEM[39788];
assign MEM[44767] = MEM[39675] + MEM[39791];
assign MEM[44768] = MEM[39676] + MEM[39717];
assign MEM[44769] = MEM[39679] + MEM[39712];
assign MEM[44770] = MEM[39680] + MEM[39780];
assign MEM[44771] = MEM[39681] + MEM[39756];
assign MEM[44772] = MEM[39682] + MEM[39801];
assign MEM[44773] = MEM[39683] + MEM[39704];
assign MEM[44774] = MEM[39684] + MEM[39708];
assign MEM[44775] = MEM[39686] + MEM[39725];
assign MEM[44776] = MEM[39687] + MEM[39758];
assign MEM[44777] = MEM[39691] + MEM[39830];
assign MEM[44778] = MEM[39692] + MEM[39732];
assign MEM[44779] = MEM[39694] + MEM[39705];
assign MEM[44780] = MEM[39697] + MEM[39815];
assign MEM[44781] = MEM[39699] + MEM[39742];
assign MEM[44782] = MEM[39700] + MEM[39883];
assign MEM[44783] = MEM[39701] + MEM[39736];
assign MEM[44784] = MEM[39702] + MEM[39724];
assign MEM[44785] = MEM[39707] + MEM[39866];
assign MEM[44786] = MEM[39709] + MEM[39718];
assign MEM[44787] = MEM[39711] + MEM[39835];
assign MEM[44788] = MEM[39713] + MEM[39739];
assign MEM[44789] = MEM[39714] + MEM[39793];
assign MEM[44790] = MEM[39719] + MEM[39753];
assign MEM[44791] = MEM[39721] + MEM[39743];
assign MEM[44792] = MEM[39722] + MEM[39821];
assign MEM[44793] = MEM[39723] + MEM[39771];
assign MEM[44794] = MEM[39728] + MEM[39737];
assign MEM[44795] = MEM[39729] + MEM[39822];
assign MEM[44796] = MEM[39730] + MEM[39785];
assign MEM[44797] = MEM[39731] + MEM[39777];
assign MEM[44798] = MEM[39733] + MEM[39757];
assign MEM[44799] = MEM[39734] + MEM[39754];
assign MEM[44800] = MEM[39735] + MEM[39797];
assign MEM[44801] = MEM[39738] + MEM[39880];
assign MEM[44802] = MEM[39740] + MEM[39890];
assign MEM[44803] = MEM[39741] + MEM[39763];
assign MEM[44804] = MEM[39744] + MEM[39798];
assign MEM[44805] = MEM[39745] + MEM[39786];
assign MEM[44806] = MEM[39746] + MEM[39810];
assign MEM[44807] = MEM[39747] + MEM[39832];
assign MEM[44808] = MEM[39748] + MEM[39767];
assign MEM[44809] = MEM[39750] + MEM[39805];
assign MEM[44810] = MEM[39751] + MEM[39770];
assign MEM[44811] = MEM[39752] + MEM[39902];
assign MEM[44812] = MEM[39755] + MEM[39870];
assign MEM[44813] = MEM[39761] + MEM[39790];
assign MEM[44814] = MEM[39762] + MEM[39808];
assign MEM[44815] = MEM[39764] + MEM[39796];
assign MEM[44816] = MEM[39765] + MEM[39827];
assign MEM[44817] = MEM[39766] + MEM[39858];
assign MEM[44818] = MEM[39768] + MEM[39823];
assign MEM[44819] = MEM[39769] + MEM[39807];
assign MEM[44820] = MEM[39772] + MEM[39960];
assign MEM[44821] = MEM[39773] + MEM[39838];
assign MEM[44822] = MEM[39774] + MEM[39789];
assign MEM[44823] = MEM[39775] + MEM[39855];
assign MEM[44824] = MEM[39776] + MEM[39897];
assign MEM[44825] = MEM[39778] + MEM[39861];
assign MEM[44826] = MEM[39779] + MEM[39837];
assign MEM[44827] = MEM[39781] + MEM[39826];
assign MEM[44828] = MEM[39782] + MEM[39851];
assign MEM[44829] = MEM[39783] + MEM[39812];
assign MEM[44830] = MEM[39784] + MEM[39872];
assign MEM[44831] = MEM[39787] + MEM[39834];
assign MEM[44832] = MEM[39792] + MEM[39828];
assign MEM[44833] = MEM[39794] + MEM[39869];
assign MEM[44834] = MEM[39799] + MEM[39811];
assign MEM[44835] = MEM[39800] + MEM[39839];
assign MEM[44836] = MEM[39802] + MEM[39840];
assign MEM[44837] = MEM[39803] + MEM[39819];
assign MEM[44838] = MEM[39804] + MEM[39895];
assign MEM[44839] = MEM[39806] + MEM[39853];
assign MEM[44840] = MEM[39809] + MEM[39977];
assign MEM[44841] = MEM[39813] + MEM[39909];
assign MEM[44842] = MEM[39814] + MEM[39891];
assign MEM[44843] = MEM[39816] + MEM[39873];
assign MEM[44844] = MEM[39817] + MEM[39871];
assign MEM[44845] = MEM[39818] + MEM[39913];
assign MEM[44846] = MEM[39820] + MEM[39863];
assign MEM[44847] = MEM[39824] + MEM[40099];
assign MEM[44848] = MEM[39825] + MEM[39995];
assign MEM[44849] = MEM[39829] + MEM[39857];
assign MEM[44850] = MEM[39831] + MEM[39947];
assign MEM[44851] = MEM[39833] + MEM[39865];
assign MEM[44852] = MEM[39841] + MEM[40069];
assign MEM[44853] = MEM[39842] + MEM[39961];
assign MEM[44854] = MEM[39843] + MEM[39915];
assign MEM[44855] = MEM[39844] + MEM[39864];
assign MEM[44856] = MEM[39845] + MEM[39914];
assign MEM[44857] = MEM[39846] + MEM[39875];
assign MEM[44858] = MEM[39847] + MEM[39963];
assign MEM[44859] = MEM[39848] + MEM[39912];
assign MEM[44860] = MEM[39849] + MEM[39881];
assign MEM[44861] = MEM[39850] + MEM[39943];
assign MEM[44862] = MEM[39852] + MEM[39899];
assign MEM[44863] = MEM[39854] + MEM[39894];
assign MEM[44864] = MEM[39856] + MEM[39916];
assign MEM[44865] = MEM[39859] + MEM[39887];
assign MEM[44866] = MEM[39860] + MEM[39922];
assign MEM[44867] = MEM[39862] + MEM[39886];
assign MEM[44868] = MEM[39867] + MEM[39901];
assign MEM[44869] = MEM[39868] + MEM[39967];
assign MEM[44870] = MEM[39874] + MEM[39879];
assign MEM[44871] = MEM[39876] + MEM[39924];
assign MEM[44872] = MEM[39877] + MEM[39970];
assign MEM[44873] = MEM[39878] + MEM[39904];
assign MEM[44874] = MEM[39882] + MEM[39964];
assign MEM[44875] = MEM[39884] + MEM[39918];
assign MEM[44876] = MEM[39885] + MEM[39923];
assign MEM[44877] = MEM[39888] + MEM[39962];
assign MEM[44878] = MEM[39889] + MEM[39898];
assign MEM[44879] = MEM[39892] + MEM[39938];
assign MEM[44880] = MEM[39893] + MEM[39944];
assign MEM[44881] = MEM[39896] + MEM[40009];
assign MEM[44882] = MEM[39900] + MEM[39930];
assign MEM[44883] = MEM[39903] + MEM[39927];
assign MEM[44884] = MEM[39905] + MEM[39979];
assign MEM[44885] = MEM[39906] + MEM[39931];
assign MEM[44886] = MEM[39907] + MEM[39950];
assign MEM[44887] = MEM[39908] + MEM[39935];
assign MEM[44888] = MEM[39910] + MEM[39949];
assign MEM[44889] = MEM[39911] + MEM[40039];
assign MEM[44890] = MEM[39917] + MEM[39934];
assign MEM[44891] = MEM[39919] + MEM[40003];
assign MEM[44892] = MEM[39920] + MEM[39953];
assign MEM[44893] = MEM[39921] + MEM[39948];
assign MEM[44894] = MEM[39925] + MEM[40051];
assign MEM[44895] = MEM[39926] + MEM[40088];
assign MEM[44896] = MEM[39928] + MEM[40052];
assign MEM[44897] = MEM[39929] + MEM[39983];
assign MEM[44898] = MEM[39932] + MEM[39975];
assign MEM[44899] = MEM[39933] + MEM[39945];
assign MEM[44900] = MEM[39936] + MEM[40071];
assign MEM[44901] = MEM[39937] + MEM[39998];
assign MEM[44902] = MEM[39939] + MEM[40008];
assign MEM[44903] = MEM[39940] + MEM[40013];
assign MEM[44904] = MEM[39941] + MEM[39958];
assign MEM[44905] = MEM[39942] + MEM[40004];
assign MEM[44906] = MEM[39946] + MEM[39966];
assign MEM[44907] = MEM[39951] + MEM[40056];
assign MEM[44908] = MEM[39952] + MEM[40010];
assign MEM[44909] = MEM[39954] + MEM[40060];
assign MEM[44910] = MEM[39955] + MEM[40054];
assign MEM[44911] = MEM[39956] + MEM[39991];
assign MEM[44912] = MEM[39957] + MEM[40082];
assign MEM[44913] = MEM[39959] + MEM[39988];
assign MEM[44914] = MEM[39965] + MEM[40103];
assign MEM[44915] = MEM[39968] + MEM[40119];
assign MEM[44916] = MEM[39969] + MEM[40091];
assign MEM[44917] = MEM[39971] + MEM[40136];
assign MEM[44918] = MEM[39972] + MEM[39996];
assign MEM[44919] = MEM[39973] + MEM[40015];
assign MEM[44920] = MEM[39974] + MEM[40025];
assign MEM[44921] = MEM[39976] + MEM[39999];
assign MEM[44922] = MEM[39978] + MEM[40017];
assign MEM[44923] = MEM[39980] + MEM[40035];
assign MEM[44924] = MEM[39981] + MEM[40043];
assign MEM[44925] = MEM[39982] + MEM[39990];
assign MEM[44926] = MEM[39984] + MEM[40094];
assign MEM[44927] = MEM[39985] + MEM[40074];
assign MEM[44928] = MEM[39986] + MEM[40041];
assign MEM[44929] = MEM[39987] + MEM[40021];
assign MEM[44930] = MEM[39989] + MEM[40005];
assign MEM[44931] = MEM[39992] + MEM[40079];
assign MEM[44932] = MEM[39993] + MEM[40040];
assign MEM[44933] = MEM[39994] + MEM[40024];
assign MEM[44934] = MEM[39997] + MEM[40102];
assign MEM[44935] = MEM[40000] + MEM[40016];
assign MEM[44936] = MEM[40001] + MEM[40037];
assign MEM[44937] = MEM[40002] + MEM[40073];
assign MEM[44938] = MEM[40006] + MEM[40028];
assign MEM[44939] = MEM[40007] + MEM[40133];
assign MEM[44940] = MEM[40011] + MEM[40062];
assign MEM[44941] = MEM[40012] + MEM[40030];
assign MEM[44942] = MEM[40014] + MEM[40061];
assign MEM[44943] = MEM[40018] + MEM[40044];
assign MEM[44944] = MEM[40019] + MEM[40034];
assign MEM[44945] = MEM[40020] + MEM[40053];
assign MEM[44946] = MEM[40022] + MEM[40195];
assign MEM[44947] = MEM[40023] + MEM[40104];
assign MEM[44948] = MEM[40026] + MEM[40108];
assign MEM[44949] = MEM[40027] + MEM[40076];
assign MEM[44950] = MEM[40029] + MEM[40095];
assign MEM[44951] = MEM[40031] + MEM[40191];
assign MEM[44952] = MEM[40032] + MEM[40065];
assign MEM[44953] = MEM[40033] + MEM[40050];
assign MEM[44954] = MEM[40036] + MEM[40057];
assign MEM[44955] = MEM[40038] + MEM[40055];
assign MEM[44956] = MEM[40042] + MEM[40072];
assign MEM[44957] = MEM[40045] + MEM[40148];
assign MEM[44958] = MEM[40046] + MEM[40161];
assign MEM[44959] = MEM[40047] + MEM[40166];
assign MEM[44960] = MEM[40048] + MEM[40132];
assign MEM[44961] = MEM[40049] + MEM[40092];
assign MEM[44962] = MEM[40058] + MEM[40090];
assign MEM[44963] = MEM[40059] + MEM[40141];
assign MEM[44964] = MEM[40063] + MEM[40131];
assign MEM[44965] = MEM[40064] + MEM[40093];
assign MEM[44966] = MEM[40066] + MEM[40145];
assign MEM[44967] = MEM[40067] + MEM[40078];
assign MEM[44968] = MEM[40068] + MEM[40077];
assign MEM[44969] = MEM[40070] + MEM[40105];
assign MEM[44970] = MEM[40075] + MEM[40110];
assign MEM[44971] = MEM[40080] + MEM[40135];
assign MEM[44972] = MEM[40081] + MEM[40142];
assign MEM[44973] = MEM[40083] + MEM[40157];
assign MEM[44974] = MEM[40084] + MEM[40112];
assign MEM[44975] = MEM[40085] + MEM[40123];
assign MEM[44976] = MEM[40086] + MEM[40134];
assign MEM[44977] = MEM[40087] + MEM[40139];
assign MEM[44978] = MEM[40089] + MEM[40098];
assign MEM[44979] = MEM[40096] + MEM[40147];
assign MEM[44980] = MEM[40097] + MEM[40163];
assign MEM[44981] = MEM[40100] + MEM[40155];
assign MEM[44982] = MEM[40101] + MEM[40238];
assign MEM[44983] = MEM[40106] + MEM[40203];
assign MEM[44984] = MEM[40107] + MEM[40175];
assign MEM[44985] = MEM[40109] + MEM[40174];
assign MEM[44986] = MEM[40111] + MEM[40122];
assign MEM[44987] = MEM[40113] + MEM[40173];
assign MEM[44988] = MEM[40114] + MEM[40187];
assign MEM[44989] = MEM[40115] + MEM[40126];
assign MEM[44990] = MEM[40116] + MEM[40162];
assign MEM[44991] = MEM[40117] + MEM[40226];
assign MEM[44992] = MEM[40118] + MEM[40170];
assign MEM[44993] = MEM[40120] + MEM[40212];
assign MEM[44994] = MEM[40121] + MEM[40206];
assign MEM[44995] = MEM[40124] + MEM[40279];
assign MEM[44996] = MEM[40125] + MEM[40278];
assign MEM[44997] = MEM[40127] + MEM[40146];
assign MEM[44998] = MEM[40128] + MEM[40159];
assign MEM[44999] = MEM[40129] + MEM[40156];
assign MEM[45000] = MEM[40130] + MEM[40198];
assign MEM[45001] = MEM[40137] + MEM[40207];
assign MEM[45002] = MEM[40138] + MEM[40168];
assign MEM[45003] = MEM[40140] + MEM[40290];
assign MEM[45004] = MEM[40143] + MEM[40154];
assign MEM[45005] = MEM[40144] + MEM[40228];
assign MEM[45006] = MEM[40149] + MEM[40172];
assign MEM[45007] = MEM[40150] + MEM[40189];
assign MEM[45008] = MEM[40151] + MEM[40185];
assign MEM[45009] = MEM[40152] + MEM[40176];
assign MEM[45010] = MEM[40153] + MEM[40180];
assign MEM[45011] = MEM[40158] + MEM[40183];
assign MEM[45012] = MEM[40160] + MEM[40231];
assign MEM[45013] = MEM[40164] + MEM[40223];
assign MEM[45014] = MEM[40165] + MEM[40202];
assign MEM[45015] = MEM[40167] + MEM[40243];
assign MEM[45016] = MEM[40169] + MEM[40235];
assign MEM[45017] = MEM[40171] + MEM[40269];
assign MEM[45018] = MEM[40177] + MEM[40297];
assign MEM[45019] = MEM[40178] + MEM[40225];
assign MEM[45020] = MEM[40179] + MEM[40186];
assign MEM[45021] = MEM[40181] + MEM[40302];
assign MEM[45022] = MEM[40182] + MEM[40210];
assign MEM[45023] = MEM[40184] + MEM[40214];
assign MEM[45024] = MEM[40188] + MEM[40342];
assign MEM[45025] = MEM[40190] + MEM[40208];
assign MEM[45026] = MEM[40192] + MEM[40254];
assign MEM[45027] = MEM[40193] + MEM[40232];
assign MEM[45028] = MEM[40194] + MEM[40250];
assign MEM[45029] = MEM[40196] + MEM[40270];
assign MEM[45030] = MEM[40197] + MEM[40343];
assign MEM[45031] = MEM[40199] + MEM[40244];
assign MEM[45032] = MEM[40200] + MEM[40241];
assign MEM[45033] = MEM[40201] + MEM[40324];
assign MEM[45034] = MEM[40204] + MEM[40236];
assign MEM[45035] = MEM[40205] + MEM[40283];
assign MEM[45036] = MEM[40209] + MEM[40303];
assign MEM[45037] = MEM[40211] + MEM[40262];
assign MEM[45038] = MEM[40213] + MEM[40272];
assign MEM[45039] = MEM[40215] + MEM[40285];
assign MEM[45040] = MEM[40216] + MEM[40305];
assign MEM[45041] = MEM[40217] + MEM[40316];
assign MEM[45042] = MEM[40218] + MEM[40334];
assign MEM[45043] = MEM[40219] + MEM[40248];
assign MEM[45044] = MEM[40220] + MEM[40280];
assign MEM[45045] = MEM[40221] + MEM[40274];
assign MEM[45046] = MEM[40222] + MEM[40230];
assign MEM[45047] = MEM[40224] + MEM[40252];
assign MEM[45048] = MEM[40227] + MEM[40255];
assign MEM[45049] = MEM[40229] + MEM[40276];
assign MEM[45050] = MEM[40233] + MEM[40357];
assign MEM[45051] = MEM[40234] + MEM[40307];
assign MEM[45052] = MEM[40237] + MEM[40359];
assign MEM[45053] = MEM[40239] + MEM[40361];
assign MEM[45054] = MEM[40240] + MEM[40286];
assign MEM[45055] = MEM[40242] + MEM[40331];
assign MEM[45056] = MEM[40245] + MEM[40256];
assign MEM[45057] = MEM[40246] + MEM[40267];
assign MEM[45058] = MEM[40247] + MEM[40332];
assign MEM[45059] = MEM[40249] + MEM[40260];
assign MEM[45060] = MEM[40251] + MEM[40288];
assign MEM[45061] = MEM[40253] + MEM[40258];
assign MEM[45062] = MEM[40257] + MEM[40309];
assign MEM[45063] = MEM[40259] + MEM[40339];
assign MEM[45064] = MEM[40261] + MEM[40304];
assign MEM[45065] = MEM[40263] + MEM[40444];
assign MEM[45066] = MEM[40264] + MEM[40292];
assign MEM[45067] = MEM[40265] + MEM[40317];
assign MEM[45068] = MEM[40266] + MEM[40373];
assign MEM[45069] = MEM[40268] + MEM[40323];
assign MEM[45070] = MEM[40271] + MEM[40296];
assign MEM[45071] = MEM[40273] + MEM[40321];
assign MEM[45072] = MEM[40275] + MEM[40406];
assign MEM[45073] = MEM[40277] + MEM[40313];
assign MEM[45074] = MEM[40281] + MEM[40358];
assign MEM[45075] = MEM[40282] + MEM[40392];
assign MEM[45076] = MEM[40284] + MEM[40350];
assign MEM[45077] = MEM[40287] + MEM[40353];
assign MEM[45078] = MEM[40289] + MEM[40318];
assign MEM[45079] = MEM[40291] + MEM[40344];
assign MEM[45080] = MEM[40293] + MEM[40301];
assign MEM[45081] = MEM[40294] + MEM[40458];
assign MEM[45082] = MEM[40295] + MEM[40356];
assign MEM[45083] = MEM[40298] + MEM[40349];
assign MEM[45084] = MEM[40299] + MEM[40364];
assign MEM[45085] = MEM[40300] + MEM[40397];
assign MEM[45086] = MEM[40306] + MEM[40430];
assign MEM[45087] = MEM[40308] + MEM[40355];
assign MEM[45088] = MEM[40310] + MEM[40385];
assign MEM[45089] = MEM[40311] + MEM[40366];
assign MEM[45090] = MEM[40312] + MEM[40354];
assign MEM[45091] = MEM[40314] + MEM[40515];
assign MEM[45092] = MEM[40315] + MEM[40328];
assign MEM[45093] = MEM[40319] + MEM[40501];
assign MEM[45094] = MEM[40320] + MEM[40413];
assign MEM[45095] = MEM[40322] + MEM[40338];
assign MEM[45096] = MEM[40325] + MEM[40340];
assign MEM[45097] = MEM[40326] + MEM[40405];
assign MEM[45098] = MEM[40327] + MEM[40386];
assign MEM[45099] = MEM[40329] + MEM[40382];
assign MEM[45100] = MEM[40330] + MEM[40363];
assign MEM[45101] = MEM[40333] + MEM[40360];
assign MEM[45102] = MEM[40335] + MEM[40370];
assign MEM[45103] = MEM[40336] + MEM[40383];
assign MEM[45104] = MEM[40337] + MEM[40400];
assign MEM[45105] = MEM[40341] + MEM[40408];
assign MEM[45106] = MEM[40345] + MEM[40391];
assign MEM[45107] = MEM[40346] + MEM[40381];
assign MEM[45108] = MEM[40347] + MEM[40431];
assign MEM[45109] = MEM[40348] + MEM[40362];
assign MEM[45110] = MEM[40351] + MEM[40371];
assign MEM[45111] = MEM[40352] + MEM[40480];
assign MEM[45112] = MEM[40365] + MEM[40390];
assign MEM[45113] = MEM[40367] + MEM[40393];
assign MEM[45114] = MEM[40368] + MEM[40487];
assign MEM[45115] = MEM[40369] + MEM[40398];
assign MEM[45116] = MEM[40372] + MEM[40426];
assign MEM[45117] = MEM[40374] + MEM[40441];
assign MEM[45118] = MEM[40375] + MEM[40502];
assign MEM[45119] = MEM[40376] + MEM[40427];
assign MEM[45120] = MEM[40377] + MEM[40476];
assign MEM[45121] = MEM[40378] + MEM[40481];
assign MEM[45122] = MEM[40379] + MEM[40409];
assign MEM[45123] = MEM[40380] + MEM[40438];
assign MEM[45124] = MEM[40384] + MEM[40451];
assign MEM[45125] = MEM[40387] + MEM[40540];
assign MEM[45126] = MEM[40388] + MEM[40442];
assign MEM[45127] = MEM[40389] + MEM[40436];
assign MEM[45128] = MEM[40394] + MEM[40421];
assign MEM[45129] = MEM[40395] + MEM[40473];
assign MEM[45130] = MEM[40396] + MEM[40454];
assign MEM[45131] = MEM[40399] + MEM[40432];
assign MEM[45132] = MEM[40401] + MEM[40460];
assign MEM[45133] = MEM[40402] + MEM[40508];
assign MEM[45134] = MEM[40403] + MEM[40477];
assign MEM[45135] = MEM[40404] + MEM[40428];
assign MEM[45136] = MEM[40407] + MEM[40498];
assign MEM[45137] = MEM[40410] + MEM[40472];
assign MEM[45138] = MEM[40411] + MEM[40435];
assign MEM[45139] = MEM[40412] + MEM[40535];
assign MEM[45140] = MEM[40414] + MEM[40450];
assign MEM[45141] = MEM[40415] + MEM[40422];
assign MEM[45142] = MEM[40416] + MEM[40546];
assign MEM[45143] = MEM[40417] + MEM[40522];
assign MEM[45144] = MEM[40418] + MEM[40440];
assign MEM[45145] = MEM[40419] + MEM[40483];
assign MEM[45146] = MEM[40420] + MEM[40459];
assign MEM[45147] = MEM[40423] + MEM[40574];
assign MEM[45148] = MEM[40424] + MEM[40489];
assign MEM[45149] = MEM[40425] + MEM[40594];
assign MEM[45150] = MEM[40429] + MEM[40494];
assign MEM[45151] = MEM[40433] + MEM[40505];
assign MEM[45152] = MEM[40434] + MEM[40488];
assign MEM[45153] = MEM[40437] + MEM[40466];
assign MEM[45154] = MEM[40439] + MEM[40539];
assign MEM[45155] = MEM[40443] + MEM[40468];
assign MEM[45156] = MEM[40445] + MEM[40520];
assign MEM[45157] = MEM[40446] + MEM[40495];
assign MEM[45158] = MEM[40447] + MEM[40514];
assign MEM[45159] = MEM[40448] + MEM[40479];
assign MEM[45160] = MEM[40449] + MEM[40563];
assign MEM[45161] = MEM[40452] + MEM[40572];
assign MEM[45162] = MEM[40453] + MEM[40475];
assign MEM[45163] = MEM[40455] + MEM[40492];
assign MEM[45164] = MEM[40456] + MEM[40478];
assign MEM[45165] = MEM[40457] + MEM[40496];
assign MEM[45166] = MEM[40461] + MEM[40557];
assign MEM[45167] = MEM[40462] + MEM[40526];
assign MEM[45168] = MEM[40463] + MEM[40573];
assign MEM[45169] = MEM[40464] + MEM[40606];
assign MEM[45170] = MEM[40465] + MEM[40504];
assign MEM[45171] = MEM[40467] + MEM[40506];
assign MEM[45172] = MEM[40469] + MEM[40513];
assign MEM[45173] = MEM[40470] + MEM[40655];
assign MEM[45174] = MEM[40471] + MEM[40527];
assign MEM[45175] = MEM[40474] + MEM[40530];
assign MEM[45176] = MEM[40482] + MEM[40584];
assign MEM[45177] = MEM[40484] + MEM[40542];
assign MEM[45178] = MEM[40485] + MEM[40552];
assign MEM[45179] = MEM[40486] + MEM[40654];
assign MEM[45180] = MEM[40490] + MEM[40518];
assign MEM[45181] = MEM[40491] + MEM[40524];
assign MEM[45182] = MEM[40493] + MEM[40556];
assign MEM[45183] = MEM[40497] + MEM[40538];
assign MEM[45184] = MEM[40499] + MEM[40532];
assign MEM[45185] = MEM[40500] + MEM[40510];
assign MEM[45186] = MEM[40503] + MEM[40549];
assign MEM[45187] = MEM[40507] + MEM[40575];
assign MEM[45188] = MEM[40509] + MEM[40568];
assign MEM[45189] = MEM[40511] + MEM[40675];
assign MEM[45190] = MEM[40512] + MEM[40634];
assign MEM[45191] = MEM[40516] + MEM[40603];
assign MEM[45192] = MEM[40517] + MEM[40636];
assign MEM[45193] = MEM[40519] + MEM[40611];
assign MEM[45194] = MEM[40521] + MEM[40646];
assign MEM[45195] = MEM[40523] + MEM[40612];
assign MEM[45196] = MEM[40525] + MEM[40599];
assign MEM[45197] = MEM[40528] + MEM[40639];
assign MEM[45198] = MEM[40529] + MEM[40562];
assign MEM[45199] = MEM[40531] + MEM[40642];
assign MEM[45200] = MEM[40533] + MEM[40613];
assign MEM[45201] = MEM[40534] + MEM[40696];
assign MEM[45202] = MEM[40536] + MEM[40580];
assign MEM[45203] = MEM[40537] + MEM[40605];
assign MEM[45204] = MEM[40541] + MEM[40601];
assign MEM[45205] = MEM[40543] + MEM[40593];
assign MEM[45206] = MEM[40544] + MEM[40566];
assign MEM[45207] = MEM[40545] + MEM[40618];
assign MEM[45208] = MEM[40547] + MEM[40592];
assign MEM[45209] = MEM[40548] + MEM[40620];
assign MEM[45210] = MEM[40550] + MEM[40564];
assign MEM[45211] = MEM[40551] + MEM[40588];
assign MEM[45212] = MEM[40553] + MEM[40641];
assign MEM[45213] = MEM[40554] + MEM[40579];
assign MEM[45214] = MEM[40555] + MEM[40669];
assign MEM[45215] = MEM[40558] + MEM[40664];
assign MEM[45216] = MEM[40559] + MEM[40598];
assign MEM[45217] = MEM[40560] + MEM[40615];
assign MEM[45218] = MEM[40561] + MEM[40650];
assign MEM[45219] = MEM[40565] + MEM[40662];
assign MEM[45220] = MEM[40567] + MEM[40581];
assign MEM[45221] = MEM[40569] + MEM[40644];
assign MEM[45222] = MEM[40570] + MEM[40623];
assign MEM[45223] = MEM[40571] + MEM[40740];
assign MEM[45224] = MEM[40576] + MEM[40625];
assign MEM[45225] = MEM[40577] + MEM[40587];
assign MEM[45226] = MEM[40578] + MEM[40652];
assign MEM[45227] = MEM[40582] + MEM[40595];
assign MEM[45228] = MEM[40583] + MEM[40600];
assign MEM[45229] = MEM[40585] + MEM[40673];
assign MEM[45230] = MEM[40586] + MEM[40619];
assign MEM[45231] = MEM[40589] + MEM[40635];
assign MEM[45232] = MEM[40590] + MEM[40729];
assign MEM[45233] = MEM[40591] + MEM[40665];
assign MEM[45234] = MEM[40596] + MEM[40656];
assign MEM[45235] = MEM[40597] + MEM[40657];
assign MEM[45236] = MEM[40602] + MEM[40626];
assign MEM[45237] = MEM[40604] + MEM[40713];
assign MEM[45238] = MEM[40607] + MEM[40629];
assign MEM[45239] = MEM[40608] + MEM[40710];
assign MEM[45240] = MEM[40609] + MEM[40697];
assign MEM[45241] = MEM[40610] + MEM[40667];
assign MEM[45242] = MEM[40614] + MEM[40632];
assign MEM[45243] = MEM[40616] + MEM[40645];
assign MEM[45244] = MEM[40617] + MEM[40622];
assign MEM[45245] = MEM[40621] + MEM[40651];
assign MEM[45246] = MEM[40624] + MEM[40700];
assign MEM[45247] = MEM[40627] + MEM[40690];
assign MEM[45248] = MEM[40628] + MEM[40707];
assign MEM[45249] = MEM[40630] + MEM[40670];
assign MEM[45250] = MEM[40631] + MEM[40774];
assign MEM[45251] = MEM[40633] + MEM[40809];
assign MEM[45252] = MEM[40637] + MEM[40771];
assign MEM[45253] = MEM[40638] + MEM[40694];
assign MEM[45254] = MEM[40640] + MEM[40743];
assign MEM[45255] = MEM[40643] + MEM[40658];
assign MEM[45256] = MEM[40647] + MEM[40704];
assign MEM[45257] = MEM[40648] + MEM[40793];
assign MEM[45258] = MEM[40649] + MEM[40679];
assign MEM[45259] = MEM[40653] + MEM[40671];
assign MEM[45260] = MEM[40659] + MEM[40734];
assign MEM[45261] = MEM[40660] + MEM[40672];
assign MEM[45262] = MEM[40661] + MEM[40686];
assign MEM[45263] = MEM[40663] + MEM[40692];
assign MEM[45264] = MEM[40666] + MEM[40685];
assign MEM[45265] = MEM[40668] + MEM[40688];
assign MEM[45266] = MEM[40674] + MEM[40687];
assign MEM[45267] = MEM[40676] + MEM[40709];
assign MEM[45268] = MEM[40677] + MEM[40744];
assign MEM[45269] = MEM[40678] + MEM[40756];
assign MEM[45270] = MEM[40680] + MEM[40750];
assign MEM[45271] = MEM[40681] + MEM[40717];
assign MEM[45272] = MEM[40682] + MEM[40770];
assign MEM[45273] = MEM[40683] + MEM[40825];
assign MEM[45274] = MEM[40684] + MEM[40701];
assign MEM[45275] = MEM[40689] + MEM[40808];
assign MEM[45276] = MEM[40691] + MEM[40714];
assign MEM[45277] = MEM[40693] + MEM[40718];
assign MEM[45278] = MEM[40695] + MEM[40781];
assign MEM[45279] = MEM[40698] + MEM[40753];
assign MEM[45280] = MEM[40699] + MEM[40769];
assign MEM[45281] = MEM[40702] + MEM[40732];
assign MEM[45282] = MEM[40703] + MEM[40780];
assign MEM[45283] = MEM[40705] + MEM[40810];
assign MEM[45284] = MEM[40706] + MEM[40777];
assign MEM[45285] = MEM[40708] + MEM[40755];
assign MEM[45286] = MEM[40711] + MEM[40846];
assign MEM[45287] = MEM[40712] + MEM[40733];
assign MEM[45288] = MEM[40715] + MEM[40776];
assign MEM[45289] = MEM[40716] + MEM[40761];
assign MEM[45290] = MEM[40719] + MEM[40775];
assign MEM[45291] = MEM[40720] + MEM[40736];
assign MEM[45292] = MEM[40721] + MEM[40739];
assign MEM[45293] = MEM[40722] + MEM[40791];
assign MEM[45294] = MEM[40723] + MEM[40786];
assign MEM[45295] = MEM[40724] + MEM[40762];
assign MEM[45296] = MEM[40725] + MEM[40843];
assign MEM[45297] = MEM[40726] + MEM[40779];
assign MEM[45298] = MEM[40727] + MEM[40768];
assign MEM[45299] = MEM[40728] + MEM[40806];
assign MEM[45300] = MEM[40730] + MEM[40867];
assign MEM[45301] = MEM[40731] + MEM[40773];
assign MEM[45302] = MEM[40735] + MEM[40752];
assign MEM[45303] = MEM[40737] + MEM[40852];
assign MEM[45304] = MEM[40738] + MEM[40751];
assign MEM[45305] = MEM[40741] + MEM[40749];
assign MEM[45306] = MEM[40742] + MEM[40747];
assign MEM[45307] = MEM[40745] + MEM[40891];
assign MEM[45308] = MEM[40746] + MEM[40767];
assign MEM[45309] = MEM[40748] + MEM[40851];
assign MEM[45310] = MEM[40754] + MEM[40866];
assign MEM[45311] = MEM[40757] + MEM[40829];
assign MEM[45312] = MEM[40758] + MEM[40948];
assign MEM[45313] = MEM[40759] + MEM[40834];
assign MEM[45314] = MEM[40760] + MEM[40820];
assign MEM[45315] = MEM[40763] + MEM[40819];
assign MEM[45316] = MEM[40764] + MEM[40822];
assign MEM[45317] = MEM[40765] + MEM[40821];
assign MEM[45318] = MEM[40766] + MEM[40835];
assign MEM[45319] = MEM[40772] + MEM[40805];
assign MEM[45320] = MEM[40778] + MEM[40782];
assign MEM[45321] = MEM[40783] + MEM[40811];
assign MEM[45322] = MEM[40784] + MEM[40848];
assign MEM[45323] = MEM[40785] + MEM[40936];
assign MEM[45324] = MEM[40787] + MEM[40906];
assign MEM[45325] = MEM[40788] + MEM[40812];
assign MEM[45326] = MEM[40789] + MEM[40799];
assign MEM[45327] = MEM[40790] + MEM[40983];
assign MEM[45328] = MEM[40792] + MEM[40838];
assign MEM[45329] = MEM[40794] + MEM[40842];
assign MEM[45330] = MEM[40795] + MEM[40861];
assign MEM[45331] = MEM[40796] + MEM[40816];
assign MEM[45332] = MEM[40797] + MEM[40850];
assign MEM[45333] = MEM[40798] + MEM[40814];
assign MEM[45334] = MEM[40800] + MEM[40944];
assign MEM[45335] = MEM[40801] + MEM[40832];
assign MEM[45336] = MEM[40802] + MEM[40919];
assign MEM[45337] = MEM[40803] + MEM[40855];
assign MEM[45338] = MEM[40804] + MEM[40823];
assign MEM[45339] = MEM[40807] + MEM[40914];
assign MEM[45340] = MEM[40813] + MEM[40856];
assign MEM[45341] = MEM[40815] + MEM[40860];
assign MEM[45342] = MEM[40817] + MEM[40836];
assign MEM[45343] = MEM[40818] + MEM[40877];
assign MEM[45344] = MEM[40824] + MEM[40870];
assign MEM[45345] = MEM[40826] + MEM[40857];
assign MEM[45346] = MEM[40827] + MEM[40954];
assign MEM[45347] = MEM[40828] + MEM[40897];
assign MEM[45348] = MEM[40830] + MEM[40879];
assign MEM[45349] = MEM[40831] + MEM[40937];
assign MEM[45350] = MEM[40833] + MEM[40885];
assign MEM[45351] = MEM[40837] + MEM[40839];
assign MEM[45352] = MEM[40840] + MEM[40847];
assign MEM[45353] = MEM[40841] + MEM[40931];
assign MEM[45354] = MEM[40844] + MEM[40868];
assign MEM[45355] = MEM[40845] + MEM[40921];
assign MEM[45356] = MEM[40849] + MEM[40872];
assign MEM[45357] = MEM[40853] + MEM[40899];
assign MEM[45358] = MEM[40854] + MEM[40910];
assign MEM[45359] = MEM[40858] + MEM[40912];
assign MEM[45360] = MEM[40859] + MEM[40947];
assign MEM[45361] = MEM[40862] + MEM[40929];
assign MEM[45362] = MEM[40863] + MEM[40928];
assign MEM[45363] = MEM[40864] + MEM[40941];
assign MEM[45364] = MEM[40865] + MEM[40971];
assign MEM[45365] = MEM[40869] + MEM[40896];
assign MEM[45366] = MEM[40871] + MEM[40907];
assign MEM[45367] = MEM[40873] + MEM[40953];
assign MEM[45368] = MEM[40874] + MEM[40883];
assign MEM[45369] = MEM[40875] + MEM[40924];
assign MEM[45370] = MEM[40876] + MEM[40913];
assign MEM[45371] = MEM[40878] + MEM[40905];
assign MEM[45372] = MEM[40880] + MEM[40915];
assign MEM[45373] = MEM[40881] + MEM[40933];
assign MEM[45374] = MEM[40882] + MEM[40930];
assign MEM[45375] = MEM[40884] + MEM[41033];
assign MEM[45376] = MEM[40886] + MEM[40898];
assign MEM[45377] = MEM[40887] + MEM[40902];
assign MEM[45378] = MEM[40888] + MEM[40949];
assign MEM[45379] = MEM[40889] + MEM[40917];
assign MEM[45380] = MEM[40890] + MEM[40909];
assign MEM[45381] = MEM[40892] + MEM[41113];
assign MEM[45382] = MEM[40893] + MEM[40908];
assign MEM[45383] = MEM[40894] + MEM[40957];
assign MEM[45384] = MEM[40895] + MEM[40911];
assign MEM[45385] = MEM[40900] + MEM[41043];
assign MEM[45386] = MEM[40901] + MEM[40963];
assign MEM[45387] = MEM[40903] + MEM[40916];
assign MEM[45388] = MEM[40904] + MEM[40945];
assign MEM[45389] = MEM[40918] + MEM[40988];
assign MEM[45390] = MEM[40920] + MEM[41014];
assign MEM[45391] = MEM[40922] + MEM[40986];
assign MEM[45392] = MEM[40923] + MEM[41018];
assign MEM[45393] = MEM[40925] + MEM[40940];
assign MEM[45394] = MEM[40926] + MEM[41001];
assign MEM[45395] = MEM[40927] + MEM[41030];
assign MEM[45396] = MEM[40932] + MEM[41013];
assign MEM[45397] = MEM[40934] + MEM[40935];
assign MEM[45398] = MEM[40938] + MEM[41012];
assign MEM[45399] = MEM[40939] + MEM[40967];
assign MEM[45400] = MEM[40942] + MEM[41011];
assign MEM[45401] = MEM[40943] + MEM[40952];
assign MEM[45402] = MEM[40946] + MEM[40997];
assign MEM[45403] = MEM[40950] + MEM[41015];
assign MEM[45404] = MEM[40951] + MEM[41026];
assign MEM[45405] = MEM[40955] + MEM[41071];
assign MEM[45406] = MEM[40956] + MEM[41004];
assign MEM[45407] = MEM[40958] + MEM[41118];
assign MEM[45408] = MEM[40959] + MEM[40998];
assign MEM[45409] = MEM[40960] + MEM[41042];
assign MEM[45410] = MEM[40961] + MEM[40999];
assign MEM[45411] = MEM[40962] + MEM[41029];
assign MEM[45412] = MEM[40964] + MEM[41022];
assign MEM[45413] = MEM[40965] + MEM[41062];
assign MEM[45414] = MEM[40966] + MEM[41049];
assign MEM[45415] = MEM[40968] + MEM[41051];
assign MEM[45416] = MEM[40969] + MEM[41076];
assign MEM[45417] = MEM[40970] + MEM[41009];
assign MEM[45418] = MEM[40972] + MEM[40994];
assign MEM[45419] = MEM[40973] + MEM[41039];
assign MEM[45420] = MEM[40974] + MEM[41020];
assign MEM[45421] = MEM[40975] + MEM[40992];
assign MEM[45422] = MEM[40976] + MEM[41091];
assign MEM[45423] = MEM[40977] + MEM[41028];
assign MEM[45424] = MEM[40978] + MEM[41044];
assign MEM[45425] = MEM[40979] + MEM[41047];
assign MEM[45426] = MEM[40980] + MEM[41046];
assign MEM[45427] = MEM[40981] + MEM[41021];
assign MEM[45428] = MEM[40982] + MEM[41006];
assign MEM[45429] = MEM[40984] + MEM[40993];
assign MEM[45430] = MEM[40985] + MEM[41082];
assign MEM[45431] = MEM[40987] + MEM[41002];
assign MEM[45432] = MEM[40989] + MEM[41010];
assign MEM[45433] = MEM[40990] + MEM[41005];
assign MEM[45434] = MEM[40991] + MEM[41085];
assign MEM[45435] = MEM[40995] + MEM[41099];
assign MEM[45436] = MEM[40996] + MEM[41053];
assign MEM[45437] = MEM[41000] + MEM[41072];
assign MEM[45438] = MEM[41003] + MEM[41132];
assign MEM[45439] = MEM[41007] + MEM[41031];
assign MEM[45440] = MEM[41008] + MEM[41035];
assign MEM[45441] = MEM[41016] + MEM[41023];
assign MEM[45442] = MEM[41017] + MEM[41052];
assign MEM[45443] = MEM[41019] + MEM[41064];
assign MEM[45444] = MEM[41024] + MEM[41200];
assign MEM[45445] = MEM[41025] + MEM[41036];
assign MEM[45446] = MEM[41027] + MEM[41125];
assign MEM[45447] = MEM[41032] + MEM[41123];
assign MEM[45448] = MEM[41034] + MEM[41079];
assign MEM[45449] = MEM[41037] + MEM[41063];
assign MEM[45450] = MEM[41038] + MEM[41103];
assign MEM[45451] = MEM[41040] + MEM[41124];
assign MEM[45452] = MEM[41041] + MEM[41068];
assign MEM[45453] = MEM[41045] + MEM[41101];
assign MEM[45454] = MEM[41048] + MEM[41104];
assign MEM[45455] = MEM[41050] + MEM[41055];
assign MEM[45456] = MEM[41054] + MEM[41127];
assign MEM[45457] = MEM[41056] + MEM[41088];
assign MEM[45458] = MEM[41057] + MEM[41168];
assign MEM[45459] = MEM[41058] + MEM[41112];
assign MEM[45460] = MEM[41059] + MEM[41179];
assign MEM[45461] = MEM[41060] + MEM[41117];
assign MEM[45462] = MEM[41061] + MEM[41070];
assign MEM[45463] = MEM[41065] + MEM[41163];
assign MEM[45464] = MEM[41066] + MEM[41135];
assign MEM[45465] = MEM[41067] + MEM[41109];
assign MEM[45466] = MEM[41069] + MEM[41145];
assign MEM[45467] = MEM[41073] + MEM[41137];
assign MEM[45468] = MEM[41074] + MEM[41139];
assign MEM[45469] = MEM[41075] + MEM[41140];
assign MEM[45470] = MEM[41077] + MEM[41108];
assign MEM[45471] = MEM[41078] + MEM[41110];
assign MEM[45472] = MEM[41080] + MEM[41193];
assign MEM[45473] = MEM[41081] + MEM[41165];
assign MEM[45474] = MEM[41083] + MEM[41150];
assign MEM[45475] = MEM[41084] + MEM[41153];
assign MEM[45476] = MEM[41086] + MEM[41185];
assign MEM[45477] = MEM[41087] + MEM[41106];
assign MEM[45478] = MEM[41089] + MEM[41151];
assign MEM[45479] = MEM[41090] + MEM[41227];
assign MEM[45480] = MEM[41092] + MEM[41144];
assign MEM[45481] = MEM[41093] + MEM[41120];
assign MEM[45482] = MEM[41094] + MEM[41166];
assign MEM[45483] = MEM[41095] + MEM[41142];
assign MEM[45484] = MEM[41096] + MEM[41190];
assign MEM[45485] = MEM[41097] + MEM[41175];
assign MEM[45486] = MEM[41098] + MEM[41171];
assign MEM[45487] = MEM[41100] + MEM[41136];
assign MEM[45488] = MEM[41102] + MEM[41128];
assign MEM[45489] = MEM[41105] + MEM[41199];
assign MEM[45490] = MEM[41107] + MEM[41138];
assign MEM[45491] = MEM[41111] + MEM[41155];
assign MEM[45492] = MEM[41114] + MEM[41198];
assign MEM[45493] = MEM[41115] + MEM[41131];
assign MEM[45494] = MEM[41116] + MEM[41211];
assign MEM[45495] = MEM[41119] + MEM[41154];
assign MEM[45496] = MEM[41121] + MEM[41226];
assign MEM[45497] = MEM[41122] + MEM[41260];
assign MEM[45498] = MEM[41126] + MEM[41241];
assign MEM[45499] = MEM[41129] + MEM[41189];
assign MEM[45500] = MEM[41130] + MEM[41158];
assign MEM[45501] = MEM[41133] + MEM[41152];
assign MEM[45502] = MEM[41134] + MEM[41255];
assign MEM[45503] = MEM[41141] + MEM[41234];
assign MEM[45504] = MEM[41143] + MEM[41164];
assign MEM[45505] = MEM[41146] + MEM[41188];
assign MEM[45506] = MEM[41147] + MEM[41184];
assign MEM[45507] = MEM[41148] + MEM[41219];
assign MEM[45508] = MEM[41149] + MEM[41287];
assign MEM[45509] = MEM[41156] + MEM[41408];
assign MEM[45510] = MEM[41157] + MEM[41186];
assign MEM[45511] = MEM[41159] + MEM[41224];
assign MEM[45512] = MEM[41160] + MEM[41206];
assign MEM[45513] = MEM[41161] + MEM[41215];
assign MEM[45514] = MEM[41162] + MEM[41174];
assign MEM[45515] = MEM[41167] + MEM[41205];
assign MEM[45516] = MEM[41169] + MEM[41347];
assign MEM[45517] = MEM[41170] + MEM[41236];
assign MEM[45518] = MEM[41172] + MEM[41240];
assign MEM[45519] = MEM[41173] + MEM[41253];
assign MEM[45520] = MEM[41176] + MEM[41196];
assign MEM[45521] = MEM[41177] + MEM[41259];
assign MEM[45522] = MEM[41178] + MEM[41309];
assign MEM[45523] = MEM[41180] + MEM[41231];
assign MEM[45524] = MEM[41181] + MEM[41248];
assign MEM[45525] = MEM[41182] + MEM[41266];
assign MEM[45526] = MEM[41183] + MEM[41222];
assign MEM[45527] = MEM[41187] + MEM[41244];
assign MEM[45528] = MEM[41191] + MEM[41237];
assign MEM[45529] = MEM[41192] + MEM[41298];
assign MEM[45530] = MEM[41194] + MEM[41218];
assign MEM[45531] = MEM[41195] + MEM[41304];
assign MEM[45532] = MEM[41197] + MEM[41369];
assign MEM[45533] = MEM[41201] + MEM[41229];
assign MEM[45534] = MEM[41202] + MEM[41225];
assign MEM[45535] = MEM[41203] + MEM[41364];
assign MEM[45536] = MEM[41204] + MEM[41334];
assign MEM[45537] = MEM[41207] + MEM[41285];
assign MEM[45538] = MEM[41208] + MEM[41272];
assign MEM[45539] = MEM[41209] + MEM[41277];
assign MEM[45540] = MEM[41210] + MEM[41302];
assign MEM[45541] = MEM[41212] + MEM[41314];
assign MEM[45542] = MEM[41213] + MEM[41278];
assign MEM[45543] = MEM[41214] + MEM[41228];
assign MEM[45544] = MEM[41216] + MEM[41335];
assign MEM[45545] = MEM[41217] + MEM[41300];
assign MEM[45546] = MEM[41220] + MEM[41449];
assign MEM[45547] = MEM[41221] + MEM[41322];
assign MEM[45548] = MEM[41223] + MEM[41292];
assign MEM[45549] = MEM[41230] + MEM[41273];
assign MEM[45550] = MEM[41232] + MEM[41286];
assign MEM[45551] = MEM[41233] + MEM[41351];
assign MEM[45552] = MEM[41235] + MEM[41284];
assign MEM[45553] = MEM[41238] + MEM[41320];
assign MEM[45554] = MEM[41239] + MEM[41261];
assign MEM[45555] = MEM[41242] + MEM[41317];
assign MEM[45556] = MEM[41243] + MEM[41289];
assign MEM[45557] = MEM[41245] + MEM[41307];
assign MEM[45558] = MEM[41246] + MEM[41276];
assign MEM[45559] = MEM[41247] + MEM[41399];
assign MEM[45560] = MEM[41249] + MEM[41305];
assign MEM[45561] = MEM[41250] + MEM[41258];
assign MEM[45562] = MEM[41251] + MEM[41339];
assign MEM[45563] = MEM[41252] + MEM[41324];
assign MEM[45564] = MEM[41254] + MEM[41271];
assign MEM[45565] = MEM[41256] + MEM[41268];
assign MEM[45566] = MEM[41257] + MEM[41341];
assign MEM[45567] = MEM[41262] + MEM[41321];
assign MEM[45568] = MEM[41263] + MEM[41374];
assign MEM[45569] = MEM[41264] + MEM[41360];
assign MEM[45570] = MEM[41265] + MEM[41340];
assign MEM[45571] = MEM[41267] + MEM[41315];
assign MEM[45572] = MEM[41269] + MEM[41410];
assign MEM[45573] = MEM[41270] + MEM[41291];
assign MEM[45574] = MEM[41274] + MEM[41332];
assign MEM[45575] = MEM[41275] + MEM[41379];
assign MEM[45576] = MEM[41279] + MEM[41362];
assign MEM[45577] = MEM[41280] + MEM[41401];
assign MEM[45578] = MEM[41281] + MEM[41367];
assign MEM[45579] = MEM[41282] + MEM[41330];
assign MEM[45580] = MEM[41283] + MEM[41333];
assign MEM[45581] = MEM[41288] + MEM[41380];
assign MEM[45582] = MEM[41290] + MEM[41311];
assign MEM[45583] = MEM[41293] + MEM[41296];
assign MEM[45584] = MEM[41294] + MEM[41346];
assign MEM[45585] = MEM[41295] + MEM[41318];
assign MEM[45586] = MEM[41297] + MEM[41303];
assign MEM[45587] = MEM[41299] + MEM[41328];
assign MEM[45588] = MEM[41301] + MEM[41471];
assign MEM[45589] = MEM[41306] + MEM[41348];
assign MEM[45590] = MEM[41308] + MEM[41352];
assign MEM[45591] = MEM[41310] + MEM[41376];
assign MEM[45592] = MEM[41312] + MEM[41378];
assign MEM[45593] = MEM[41313] + MEM[41342];
assign MEM[45594] = MEM[41316] + MEM[41363];
assign MEM[45595] = MEM[41319] + MEM[41323];
assign MEM[45596] = MEM[41325] + MEM[41358];
assign MEM[45597] = MEM[41326] + MEM[41361];
assign MEM[45598] = MEM[41327] + MEM[41373];
assign MEM[45599] = MEM[41329] + MEM[41343];
assign MEM[45600] = MEM[41331] + MEM[41553];
assign MEM[45601] = MEM[41336] + MEM[41404];
assign MEM[45602] = MEM[41337] + MEM[41395];
assign MEM[45603] = MEM[41338] + MEM[41393];
assign MEM[45604] = MEM[41344] + MEM[41394];
assign MEM[45605] = MEM[41345] + MEM[41403];
assign MEM[45606] = MEM[41349] + MEM[41494];
assign MEM[45607] = MEM[41350] + MEM[41459];
assign MEM[45608] = MEM[41353] + MEM[41411];
assign MEM[45609] = MEM[41354] + MEM[41406];
assign MEM[45610] = MEM[41355] + MEM[41402];
assign MEM[45611] = MEM[41356] + MEM[41412];
assign MEM[45612] = MEM[41357] + MEM[41381];
assign MEM[45613] = MEM[41359] + MEM[41372];
assign MEM[45614] = MEM[41365] + MEM[41405];
assign MEM[45615] = MEM[41366] + MEM[41433];
assign MEM[45616] = MEM[41368] + MEM[41429];
assign MEM[45617] = MEM[41370] + MEM[41375];
assign MEM[45618] = MEM[41371] + MEM[41398];
assign MEM[45619] = MEM[41377] + MEM[41436];
assign MEM[45620] = MEM[41382] + MEM[41397];
assign MEM[45621] = MEM[41383] + MEM[41389];
assign MEM[45622] = MEM[41384] + MEM[41450];
assign MEM[45623] = MEM[41385] + MEM[41570];
assign MEM[45624] = MEM[41386] + MEM[41424];
assign MEM[45625] = MEM[41387] + MEM[41523];
assign MEM[45626] = MEM[41388] + MEM[41416];
assign MEM[45627] = MEM[41390] + MEM[41477];
assign MEM[45628] = MEM[41391] + MEM[41407];
assign MEM[45629] = MEM[41392] + MEM[41455];
assign MEM[45630] = MEM[41396] + MEM[41500];
assign MEM[45631] = MEM[41400] + MEM[41479];
assign MEM[45632] = MEM[41409] + MEM[41492];
assign MEM[45633] = MEM[41413] + MEM[41473];
assign MEM[45634] = MEM[41414] + MEM[41439];
assign MEM[45635] = MEM[41415] + MEM[41465];
assign MEM[45636] = MEM[41417] + MEM[41493];
assign MEM[45637] = MEM[41418] + MEM[41451];
assign MEM[45638] = MEM[41419] + MEM[41448];
assign MEM[45639] = MEM[41420] + MEM[41454];
assign MEM[45640] = MEM[41421] + MEM[41544];
assign MEM[45641] = MEM[41422] + MEM[41456];
assign MEM[45642] = MEM[41423] + MEM[41503];
assign MEM[45643] = MEM[41425] + MEM[41514];
assign MEM[45644] = MEM[41426] + MEM[41434];
assign MEM[45645] = MEM[41427] + MEM[41587];
assign MEM[45646] = MEM[41428] + MEM[41472];
assign MEM[45647] = MEM[41430] + MEM[41464];
assign MEM[45648] = MEM[41431] + MEM[41476];
assign MEM[45649] = MEM[41432] + MEM[41469];
assign MEM[45650] = MEM[41435] + MEM[41507];
assign MEM[45651] = MEM[41437] + MEM[41491];
assign MEM[45652] = MEM[41438] + MEM[41541];
assign MEM[45653] = MEM[41440] + MEM[41481];
assign MEM[45654] = MEM[41441] + MEM[41555];
assign MEM[45655] = MEM[41442] + MEM[41486];
assign MEM[45656] = MEM[41443] + MEM[41485];
assign MEM[45657] = MEM[41444] + MEM[41499];
assign MEM[45658] = MEM[41445] + MEM[41457];
assign MEM[45659] = MEM[41446] + MEM[41556];
assign MEM[45660] = MEM[41447] + MEM[41489];
assign MEM[45661] = MEM[41452] + MEM[41590];
assign MEM[45662] = MEM[41453] + MEM[41480];
assign MEM[45663] = MEM[41458] + MEM[41549];
assign MEM[45664] = MEM[41460] + MEM[41483];
assign MEM[45665] = MEM[41461] + MEM[41501];
assign MEM[45666] = MEM[41462] + MEM[41552];
assign MEM[45667] = MEM[41463] + MEM[41535];
assign MEM[45668] = MEM[41466] + MEM[41558];
assign MEM[45669] = MEM[41467] + MEM[41608];
assign MEM[45670] = MEM[41468] + MEM[41513];
assign MEM[45671] = MEM[41470] + MEM[41561];
assign MEM[45672] = MEM[41474] + MEM[41592];
assign MEM[45673] = MEM[41475] + MEM[41502];
assign MEM[45674] = MEM[41478] + MEM[41521];
assign MEM[45675] = MEM[41482] + MEM[41528];
assign MEM[45676] = MEM[41484] + MEM[41551];
assign MEM[45677] = MEM[41487] + MEM[41571];
assign MEM[45678] = MEM[41488] + MEM[41554];
assign MEM[45679] = MEM[41490] + MEM[41498];
assign MEM[45680] = MEM[41495] + MEM[41529];
assign MEM[45681] = MEM[41496] + MEM[41542];
assign MEM[45682] = MEM[41497] + MEM[41602];
assign MEM[45683] = MEM[41504] + MEM[41548];
assign MEM[45684] = MEM[41505] + MEM[41668];
assign MEM[45685] = MEM[41506] + MEM[41533];
assign MEM[45686] = MEM[41508] + MEM[41560];
assign MEM[45687] = MEM[41509] + MEM[41586];
assign MEM[45688] = MEM[41510] + MEM[41530];
assign MEM[45689] = MEM[41511] + MEM[41578];
assign MEM[45690] = MEM[41512] + MEM[41617];
assign MEM[45691] = MEM[41515] + MEM[41580];
assign MEM[45692] = MEM[41516] + MEM[41575];
assign MEM[45693] = MEM[41517] + MEM[41564];
assign MEM[45694] = MEM[41518] + MEM[41582];
assign MEM[45695] = MEM[41519] + MEM[41537];
assign MEM[45696] = MEM[41520] + MEM[41543];
assign MEM[45697] = MEM[41522] + MEM[41594];
assign MEM[45698] = MEM[41524] + MEM[41531];
assign MEM[45699] = MEM[41525] + MEM[41550];
assign MEM[45700] = MEM[41526] + MEM[41599];
assign MEM[45701] = MEM[41527] + MEM[41696];
assign MEM[45702] = MEM[41532] + MEM[41666];
assign MEM[45703] = MEM[41534] + MEM[41540];
assign MEM[45704] = MEM[41536] + MEM[41607];
assign MEM[45705] = MEM[41538] + MEM[41670];
assign MEM[45706] = MEM[41539] + MEM[41632];
assign MEM[45707] = MEM[41545] + MEM[41569];
assign MEM[45708] = MEM[41546] + MEM[41579];
assign MEM[45709] = MEM[41547] + MEM[41597];
assign MEM[45710] = MEM[41557] + MEM[41658];
assign MEM[45711] = MEM[41559] + MEM[41581];
assign MEM[45712] = MEM[41562] + MEM[41630];
assign MEM[45713] = MEM[41563] + MEM[41595];
assign MEM[45714] = MEM[41565] + MEM[41605];
assign MEM[45715] = MEM[41566] + MEM[41709];
assign MEM[45716] = MEM[41567] + MEM[41643];
assign MEM[45717] = MEM[41568] + MEM[41652];
assign MEM[45718] = MEM[41572] + MEM[41621];
assign MEM[45719] = MEM[41573] + MEM[41619];
assign MEM[45720] = MEM[41574] + MEM[41667];
assign MEM[45721] = MEM[41576] + MEM[41690];
assign MEM[45722] = MEM[41577] + MEM[41604];
assign MEM[45723] = MEM[41583] + MEM[41656];
assign MEM[45724] = MEM[41584] + MEM[41596];
assign MEM[45725] = MEM[41585] + MEM[41612];
assign MEM[45726] = MEM[41588] + MEM[41625];
assign MEM[45727] = MEM[41589] + MEM[41620];
assign MEM[45728] = MEM[41591] + MEM[41637];
assign MEM[45729] = MEM[41593] + MEM[41628];
assign MEM[45730] = MEM[41598] + MEM[41650];
assign MEM[45731] = MEM[41600] + MEM[41653];
assign MEM[45732] = MEM[41601] + MEM[41623];
assign MEM[45733] = MEM[41603] + MEM[41648];
assign MEM[45734] = MEM[41606] + MEM[41755];
assign MEM[45735] = MEM[41609] + MEM[41665];
assign MEM[45736] = MEM[41610] + MEM[41624];
assign MEM[45737] = MEM[41611] + MEM[41683];
assign MEM[45738] = MEM[41613] + MEM[41669];
assign MEM[45739] = MEM[41614] + MEM[41635];
assign MEM[45740] = MEM[41615] + MEM[41645];
assign MEM[45741] = MEM[41616] + MEM[41717];
assign MEM[45742] = MEM[41618] + MEM[41641];
assign MEM[45743] = MEM[41622] + MEM[41646];
assign MEM[45744] = MEM[41626] + MEM[41734];
assign MEM[45745] = MEM[41627] + MEM[41675];
assign MEM[45746] = MEM[41629] + MEM[41662];
assign MEM[45747] = MEM[41631] + MEM[41758];
assign MEM[45748] = MEM[41633] + MEM[41716];
assign MEM[45749] = MEM[41634] + MEM[41706];
assign MEM[45750] = MEM[41636] + MEM[41663];
assign MEM[45751] = MEM[41638] + MEM[41655];
assign MEM[45752] = MEM[41639] + MEM[41700];
assign MEM[45753] = MEM[41640] + MEM[41679];
assign MEM[45754] = MEM[41642] + MEM[41725];
assign MEM[45755] = MEM[41644] + MEM[41699];
assign MEM[45756] = MEM[41647] + MEM[41752];
assign MEM[45757] = MEM[41649] + MEM[41686];
assign MEM[45758] = MEM[41651] + MEM[41714];
assign MEM[45759] = MEM[41654] + MEM[41701];
assign MEM[45760] = MEM[41657] + MEM[41676];
assign MEM[45761] = MEM[41659] + MEM[41800];
assign MEM[45762] = MEM[41660] + MEM[41689];
assign MEM[45763] = MEM[41661] + MEM[41692];
assign MEM[45764] = MEM[41664] + MEM[41705];
assign MEM[45765] = MEM[41671] + MEM[41735];
assign MEM[45766] = MEM[41672] + MEM[41768];
assign MEM[45767] = MEM[41673] + MEM[41703];
assign MEM[45768] = MEM[41674] + MEM[41708];
assign MEM[45769] = MEM[41677] + MEM[41722];
assign MEM[45770] = MEM[41678] + MEM[41743];
assign MEM[45771] = MEM[41680] + MEM[41694];
assign MEM[45772] = MEM[41681] + MEM[41781];
assign MEM[45773] = MEM[41682] + MEM[41739];
assign MEM[45774] = MEM[41684] + MEM[41825];
assign MEM[45775] = MEM[41685] + MEM[41778];
assign MEM[45776] = MEM[41687] + MEM[41729];
assign MEM[45777] = MEM[41688] + MEM[41759];
assign MEM[45778] = MEM[41691] + MEM[41738];
assign MEM[45779] = MEM[41693] + MEM[41815];
assign MEM[45780] = MEM[41695] + MEM[41711];
assign MEM[45781] = MEM[41697] + MEM[41732];
assign MEM[45782] = MEM[41698] + MEM[41720];
assign MEM[45783] = MEM[41702] + MEM[41762];
assign MEM[45784] = MEM[41704] + MEM[41715];
assign MEM[45785] = MEM[41707] + MEM[41749];
assign MEM[45786] = MEM[41710] + MEM[41777];
assign MEM[45787] = MEM[41712] + MEM[41783];
assign MEM[45788] = MEM[41713] + MEM[41748];
assign MEM[45789] = MEM[41718] + MEM[41797];
assign MEM[45790] = MEM[41719] + MEM[41727];
assign MEM[45791] = MEM[41721] + MEM[41782];
assign MEM[45792] = MEM[41723] + MEM[41793];
assign MEM[45793] = MEM[41724] + MEM[41751];
assign MEM[45794] = MEM[41726] + MEM[41746];
assign MEM[45795] = MEM[41728] + MEM[41831];
assign MEM[45796] = MEM[41730] + MEM[41836];
assign MEM[45797] = MEM[41731] + MEM[41747];
assign MEM[45798] = MEM[41733] + MEM[41820];
assign MEM[45799] = MEM[41736] + MEM[41756];
assign MEM[45800] = MEM[41737] + MEM[41842];
assign MEM[45801] = MEM[41740] + MEM[41796];
assign MEM[45802] = MEM[41741] + MEM[41829];
assign MEM[45803] = MEM[41742] + MEM[41767];
assign MEM[45804] = MEM[41744] + MEM[41772];
assign MEM[45805] = MEM[41745] + MEM[41810];
assign MEM[45806] = MEM[41750] + MEM[41928];
assign MEM[45807] = MEM[41753] + MEM[41787];
assign MEM[45808] = MEM[41754] + MEM[41846];
assign MEM[45809] = MEM[41757] + MEM[41804];
assign MEM[45810] = MEM[41760] + MEM[41812];
assign MEM[45811] = MEM[41761] + MEM[41845];
assign MEM[45812] = MEM[41763] + MEM[41801];
assign MEM[45813] = MEM[41764] + MEM[41803];
assign MEM[45814] = MEM[41765] + MEM[41837];
assign MEM[45815] = MEM[41766] + MEM[41814];
assign MEM[45816] = MEM[41769] + MEM[41895];
assign MEM[45817] = MEM[41770] + MEM[41865];
assign MEM[45818] = MEM[41771] + MEM[41788];
assign MEM[45819] = MEM[41773] + MEM[41840];
assign MEM[45820] = MEM[41774] + MEM[41798];
assign MEM[45821] = MEM[41775] + MEM[41802];
assign MEM[45822] = MEM[41776] + MEM[41860];
assign MEM[45823] = MEM[41779] + MEM[41806];
assign MEM[45824] = MEM[41780] + MEM[41816];
assign MEM[45825] = MEM[41784] + MEM[41857];
assign MEM[45826] = MEM[41785] + MEM[41869];
assign MEM[45827] = MEM[41786] + MEM[41826];
assign MEM[45828] = MEM[41789] + MEM[41910];
assign MEM[45829] = MEM[41790] + MEM[41834];
assign MEM[45830] = MEM[41791] + MEM[41883];
assign MEM[45831] = MEM[41792] + MEM[41823];
assign MEM[45832] = MEM[41794] + MEM[41851];
assign MEM[45833] = MEM[41795] + MEM[41917];
assign MEM[45834] = MEM[41799] + MEM[41841];
assign MEM[45835] = MEM[41805] + MEM[41830];
assign MEM[45836] = MEM[41807] + MEM[41891];
assign MEM[45837] = MEM[41808] + MEM[41849];
assign MEM[45838] = MEM[41809] + MEM[41916];
assign MEM[45839] = MEM[41811] + MEM[41922];
assign MEM[45840] = MEM[41813] + MEM[41874];
assign MEM[45841] = MEM[41817] + MEM[41856];
assign MEM[45842] = MEM[41818] + MEM[41906];
assign MEM[45843] = MEM[41819] + MEM[41934];
assign MEM[45844] = MEM[41821] + MEM[41832];
assign MEM[45845] = MEM[41822] + MEM[41926];
assign MEM[45846] = MEM[41824] + MEM[41838];
assign MEM[45847] = MEM[41827] + MEM[41875];
assign MEM[45848] = MEM[41828] + MEM[41939];
assign MEM[45849] = MEM[41833] + MEM[41893];
assign MEM[45850] = MEM[41835] + MEM[41959];
assign MEM[45851] = MEM[41839] + MEM[41848];
assign MEM[45852] = MEM[41843] + MEM[41876];
assign MEM[45853] = MEM[41844] + MEM[41923];
assign MEM[45854] = MEM[41847] + MEM[41861];
assign MEM[45855] = MEM[41850] + MEM[41900];
assign MEM[45856] = MEM[41852] + MEM[41932];
assign MEM[45857] = MEM[41853] + MEM[41911];
assign MEM[45858] = MEM[41854] + MEM[41889];
assign MEM[45859] = MEM[41855] + MEM[41892];
assign MEM[45860] = MEM[41858] + MEM[41940];
assign MEM[45861] = MEM[41859] + MEM[41909];
assign MEM[45862] = MEM[41862] + MEM[41927];
assign MEM[45863] = MEM[41863] + MEM[41930];
assign MEM[45864] = MEM[41864] + MEM[41956];
assign MEM[45865] = MEM[41866] + MEM[41897];
assign MEM[45866] = MEM[41867] + MEM[41888];
assign MEM[45867] = MEM[41868] + MEM[41899];
assign MEM[45868] = MEM[41870] + MEM[41907];
assign MEM[45869] = MEM[41871] + MEM[41965];
assign MEM[45870] = MEM[41872] + MEM[41898];
assign MEM[45871] = MEM[41873] + MEM[41938];
assign MEM[45872] = MEM[41877] + MEM[41920];
assign MEM[45873] = MEM[41878] + MEM[41894];
assign MEM[45874] = MEM[41879] + MEM[41915];
assign MEM[45875] = MEM[41880] + MEM[41937];
assign MEM[45876] = MEM[41881] + MEM[41960];
assign MEM[45877] = MEM[41882] + MEM[41981];
assign MEM[45878] = MEM[41884] + MEM[42011];
assign MEM[45879] = MEM[41885] + MEM[41952];
assign MEM[45880] = MEM[41886] + MEM[41941];
assign MEM[45881] = MEM[41887] + MEM[41993];
assign MEM[45882] = MEM[41890] + MEM[41924];
assign MEM[45883] = MEM[41896] + MEM[41977];
assign MEM[45884] = MEM[41901] + MEM[41948];
assign MEM[45885] = MEM[41902] + MEM[41970];
assign MEM[45886] = MEM[41903] + MEM[41951];
assign MEM[45887] = MEM[41904] + MEM[41996];
assign MEM[45888] = MEM[41905] + MEM[42036];
assign MEM[45889] = MEM[41908] + MEM[41999];
assign MEM[45890] = MEM[41912] + MEM[42007];
assign MEM[45891] = MEM[41913] + MEM[41936];
assign MEM[45892] = MEM[41914] + MEM[42010];
assign MEM[45893] = MEM[41918] + MEM[41986];
assign MEM[45894] = MEM[41919] + MEM[41943];
assign MEM[45895] = MEM[41921] + MEM[41955];
assign MEM[45896] = MEM[41925] + MEM[41961];
assign MEM[45897] = MEM[41929] + MEM[41972];
assign MEM[45898] = MEM[41931] + MEM[41958];
assign MEM[45899] = MEM[41933] + MEM[41984];
assign MEM[45900] = MEM[41935] + MEM[41953];
assign MEM[45901] = MEM[41942] + MEM[41947];
assign MEM[45902] = MEM[41944] + MEM[42027];
assign MEM[45903] = MEM[41945] + MEM[42066];
assign MEM[45904] = MEM[41946] + MEM[42044];
assign MEM[45905] = MEM[41949] + MEM[42032];
assign MEM[45906] = MEM[41950] + MEM[41982];
assign MEM[45907] = MEM[41954] + MEM[42015];
assign MEM[45908] = MEM[41957] + MEM[42019];
assign MEM[45909] = MEM[41962] + MEM[42041];
assign MEM[45910] = MEM[41963] + MEM[41990];
assign MEM[45911] = MEM[41964] + MEM[42034];
assign MEM[45912] = MEM[41966] + MEM[42004];
assign MEM[45913] = MEM[41967] + MEM[42076];
assign MEM[45914] = MEM[41968] + MEM[42046];
assign MEM[45915] = MEM[41969] + MEM[42033];
assign MEM[45916] = MEM[41971] + MEM[42029];
assign MEM[45917] = MEM[41973] + MEM[42047];
assign MEM[45918] = MEM[41974] + MEM[42050];
assign MEM[45919] = MEM[41975] + MEM[42085];
assign MEM[45920] = MEM[41976] + MEM[42071];
assign MEM[45921] = MEM[41978] + MEM[42003];
assign MEM[45922] = MEM[41979] + MEM[42035];
assign MEM[45923] = MEM[41980] + MEM[42049];
assign MEM[45924] = MEM[41983] + MEM[42177];
assign MEM[45925] = MEM[41985] + MEM[41998];
assign MEM[45926] = MEM[41987] + MEM[42078];
assign MEM[45927] = MEM[41988] + MEM[42054];
assign MEM[45928] = MEM[41989] + MEM[42026];
assign MEM[45929] = MEM[41991] + MEM[42059];
assign MEM[45930] = MEM[41992] + MEM[42001];
assign MEM[45931] = MEM[41994] + MEM[42112];
assign MEM[45932] = MEM[41995] + MEM[42028];
assign MEM[45933] = MEM[41997] + MEM[42022];
assign MEM[45934] = MEM[42000] + MEM[42018];
assign MEM[45935] = MEM[42002] + MEM[42043];
assign MEM[45936] = MEM[42005] + MEM[42065];
assign MEM[45937] = MEM[42006] + MEM[42095];
assign MEM[45938] = MEM[42008] + MEM[42072];
assign MEM[45939] = MEM[42009] + MEM[42081];
assign MEM[45940] = MEM[42012] + MEM[42070];
assign MEM[45941] = MEM[42013] + MEM[42060];
assign MEM[45942] = MEM[42014] + MEM[42058];
assign MEM[45943] = MEM[42016] + MEM[42073];
assign MEM[45944] = MEM[42017] + MEM[42038];
assign MEM[45945] = MEM[42020] + MEM[42057];
assign MEM[45946] = MEM[42021] + MEM[42053];
assign MEM[45947] = MEM[42023] + MEM[42111];
assign MEM[45948] = MEM[42024] + MEM[42099];
assign MEM[45949] = MEM[42025] + MEM[42101];
assign MEM[45950] = MEM[42030] + MEM[42105];
assign MEM[45951] = MEM[42031] + MEM[42216];
assign MEM[45952] = MEM[42037] + MEM[42109];
assign MEM[45953] = MEM[42039] + MEM[42087];
assign MEM[45954] = MEM[42040] + MEM[42184];
assign MEM[45955] = MEM[42042] + MEM[42074];
assign MEM[45956] = MEM[42045] + MEM[42132];
assign MEM[45957] = MEM[42048] + MEM[42090];
assign MEM[45958] = MEM[42051] + MEM[42110];
assign MEM[45959] = MEM[42052] + MEM[42098];
assign MEM[45960] = MEM[42055] + MEM[42106];
assign MEM[45961] = MEM[42056] + MEM[42116];
assign MEM[45962] = MEM[42061] + MEM[42083];
assign MEM[45963] = MEM[42062] + MEM[42104];
assign MEM[45964] = MEM[42063] + MEM[42147];
assign MEM[45965] = MEM[42064] + MEM[42137];
assign MEM[45966] = MEM[42067] + MEM[42173];
assign MEM[45967] = MEM[42068] + MEM[42118];
assign MEM[45968] = MEM[42069] + MEM[42080];
assign MEM[45969] = MEM[42075] + MEM[42121];
assign MEM[45970] = MEM[42077] + MEM[42094];
assign MEM[45971] = MEM[42079] + MEM[42162];
assign MEM[45972] = MEM[42082] + MEM[42181];
assign MEM[45973] = MEM[42084] + MEM[42113];
assign MEM[45974] = MEM[42086] + MEM[42185];
assign MEM[45975] = MEM[42088] + MEM[42103];
assign MEM[45976] = MEM[42089] + MEM[42222];
assign MEM[45977] = MEM[42091] + MEM[42126];
assign MEM[45978] = MEM[42092] + MEM[42148];
assign MEM[45979] = MEM[42093] + MEM[42125];
assign MEM[45980] = MEM[42096] + MEM[42142];
assign MEM[45981] = MEM[42097] + MEM[42169];
assign MEM[45982] = MEM[42100] + MEM[42127];
assign MEM[45983] = MEM[42102] + MEM[42152];
assign MEM[45984] = MEM[42107] + MEM[42163];
assign MEM[45985] = MEM[42108] + MEM[42200];
assign MEM[45986] = MEM[42114] + MEM[42122];
assign MEM[45987] = MEM[42115] + MEM[42194];
assign MEM[45988] = MEM[42117] + MEM[42154];
assign MEM[45989] = MEM[42119] + MEM[42139];
assign MEM[45990] = MEM[42120] + MEM[42191];
assign MEM[45991] = MEM[42123] + MEM[42171];
assign MEM[45992] = MEM[42124] + MEM[42219];
assign MEM[45993] = MEM[42128] + MEM[42160];
assign MEM[45994] = MEM[42129] + MEM[42175];
assign MEM[45995] = MEM[42130] + MEM[42141];
assign MEM[45996] = MEM[42131] + MEM[42252];
assign MEM[45997] = MEM[42133] + MEM[42221];
assign MEM[45998] = MEM[42134] + MEM[42284];
assign MEM[45999] = MEM[42135] + MEM[42165];
assign MEM[46000] = MEM[42136] + MEM[42270];
assign MEM[46001] = MEM[42138] + MEM[42187];
assign MEM[46002] = MEM[42140] + MEM[42214];
assign MEM[46003] = MEM[42143] + MEM[42182];
assign MEM[46004] = MEM[42144] + MEM[42271];
assign MEM[46005] = MEM[42145] + MEM[42201];
assign MEM[46006] = MEM[42146] + MEM[42196];
assign MEM[46007] = MEM[42149] + MEM[42193];
assign MEM[46008] = MEM[42150] + MEM[42192];
assign MEM[46009] = MEM[42151] + MEM[42203];
assign MEM[46010] = MEM[42153] + MEM[42238];
assign MEM[46011] = MEM[42155] + MEM[42178];
assign MEM[46012] = MEM[42156] + MEM[42236];
assign MEM[46013] = MEM[42157] + MEM[42189];
assign MEM[46014] = MEM[42158] + MEM[42241];
assign MEM[46015] = MEM[42159] + MEM[42230];
assign MEM[46016] = MEM[42161] + MEM[42218];
assign MEM[46017] = MEM[42164] + MEM[42199];
assign MEM[46018] = MEM[42166] + MEM[42195];
assign MEM[46019] = MEM[42167] + MEM[42211];
assign MEM[46020] = MEM[42168] + MEM[42179];
assign MEM[46021] = MEM[42170] + MEM[42248];
assign MEM[46022] = MEM[42172] + MEM[42225];
assign MEM[46023] = MEM[42174] + MEM[42316];
assign MEM[46024] = MEM[42176] + MEM[42240];
assign MEM[46025] = MEM[42180] + MEM[42204];
assign MEM[46026] = MEM[42183] + MEM[42229];
assign MEM[46027] = MEM[42186] + MEM[42242];
assign MEM[46028] = MEM[42188] + MEM[42268];
assign MEM[46029] = MEM[42190] + MEM[42250];
assign MEM[46030] = MEM[42197] + MEM[42224];
assign MEM[46031] = MEM[42198] + MEM[42265];
assign MEM[46032] = MEM[42202] + MEM[42303];
assign MEM[46033] = MEM[42205] + MEM[42319];
assign MEM[46034] = MEM[42206] + MEM[42273];
assign MEM[46035] = MEM[42207] + MEM[42239];
assign MEM[46036] = MEM[42208] + MEM[42259];
assign MEM[46037] = MEM[42209] + MEM[42278];
assign MEM[46038] = MEM[42210] + MEM[42261];
assign MEM[46039] = MEM[42212] + MEM[42282];
assign MEM[46040] = MEM[42213] + MEM[42285];
assign MEM[46041] = MEM[42215] + MEM[42256];
assign MEM[46042] = MEM[42217] + MEM[42276];
assign MEM[46043] = MEM[42220] + MEM[42311];
assign MEM[46044] = MEM[42223] + MEM[42292];
assign MEM[46045] = MEM[42226] + MEM[42266];
assign MEM[46046] = MEM[42227] + MEM[42297];
assign MEM[46047] = MEM[42228] + MEM[42300];
assign MEM[46048] = MEM[42231] + MEM[42337];
assign MEM[46049] = MEM[42232] + MEM[42244];
assign MEM[46050] = MEM[42233] + MEM[42260];
assign MEM[46051] = MEM[42234] + MEM[42269];
assign MEM[46052] = MEM[42235] + MEM[42247];
assign MEM[46053] = MEM[42237] + MEM[42310];
assign MEM[46054] = MEM[42243] + MEM[42264];
assign MEM[46055] = MEM[42245] + MEM[42408];
assign MEM[46056] = MEM[42246] + MEM[42291];
assign MEM[46057] = MEM[42249] + MEM[42263];
assign MEM[46058] = MEM[42251] + MEM[42348];
assign MEM[46059] = MEM[42253] + MEM[42386];
assign MEM[46060] = MEM[42254] + MEM[42288];
assign MEM[46061] = MEM[42255] + MEM[42346];
assign MEM[46062] = MEM[42257] + MEM[42350];
assign MEM[46063] = MEM[42258] + MEM[42344];
assign MEM[46064] = MEM[42262] + MEM[42286];
assign MEM[46065] = MEM[42267] + MEM[42349];
assign MEM[46066] = MEM[42272] + MEM[42356];
assign MEM[46067] = MEM[42274] + MEM[42425];
assign MEM[46068] = MEM[42275] + MEM[42336];
assign MEM[46069] = MEM[42277] + MEM[42294];
assign MEM[46070] = MEM[42279] + MEM[42334];
assign MEM[46071] = MEM[42280] + MEM[42393];
assign MEM[46072] = MEM[42281] + MEM[42382];
assign MEM[46073] = MEM[42283] + MEM[42345];
assign MEM[46074] = MEM[42287] + MEM[42374];
assign MEM[46075] = MEM[42289] + MEM[42329];
assign MEM[46076] = MEM[42290] + MEM[42308];
assign MEM[46077] = MEM[42293] + MEM[42335];
assign MEM[46078] = MEM[42295] + MEM[42362];
assign MEM[46079] = MEM[42296] + MEM[42324];
assign MEM[46080] = MEM[42298] + MEM[42342];
assign MEM[46081] = MEM[42299] + MEM[42368];
assign MEM[46082] = MEM[42301] + MEM[42445];
assign MEM[46083] = MEM[42302] + MEM[42419];
assign MEM[46084] = MEM[42304] + MEM[42347];
assign MEM[46085] = MEM[42305] + MEM[42387];
assign MEM[46086] = MEM[42306] + MEM[42352];
assign MEM[46087] = MEM[42307] + MEM[42326];
assign MEM[46088] = MEM[42309] + MEM[42372];
assign MEM[46089] = MEM[42312] + MEM[42379];
assign MEM[46090] = MEM[42313] + MEM[42460];
assign MEM[46091] = MEM[42314] + MEM[42358];
assign MEM[46092] = MEM[42315] + MEM[42365];
assign MEM[46093] = MEM[42317] + MEM[42354];
assign MEM[46094] = MEM[42318] + MEM[42414];
assign MEM[46095] = MEM[42320] + MEM[42366];
assign MEM[46096] = MEM[42321] + MEM[42385];
assign MEM[46097] = MEM[42322] + MEM[42412];
assign MEM[46098] = MEM[42323] + MEM[42369];
assign MEM[46099] = MEM[42325] + MEM[42351];
assign MEM[46100] = MEM[42327] + MEM[42396];
assign MEM[46101] = MEM[42328] + MEM[42364];
assign MEM[46102] = MEM[42330] + MEM[42418];
assign MEM[46103] = MEM[42331] + MEM[42429];
assign MEM[46104] = MEM[42332] + MEM[42373];
assign MEM[46105] = MEM[42333] + MEM[42367];
assign MEM[46106] = MEM[42338] + MEM[42391];
assign MEM[46107] = MEM[42339] + MEM[42437];
assign MEM[46108] = MEM[42340] + MEM[42376];
assign MEM[46109] = MEM[42341] + MEM[42375];
assign MEM[46110] = MEM[42343] + MEM[42381];
assign MEM[46111] = MEM[42353] + MEM[42469];
assign MEM[46112] = MEM[42355] + MEM[42433];
assign MEM[46113] = MEM[42357] + MEM[42404];
assign MEM[46114] = MEM[42359] + MEM[42405];
assign MEM[46115] = MEM[42360] + MEM[42432];
assign MEM[46116] = MEM[42361] + MEM[42383];
assign MEM[46117] = MEM[42363] + MEM[42409];
assign MEM[46118] = MEM[42370] + MEM[42454];
assign MEM[46119] = MEM[42371] + MEM[42421];
assign MEM[46120] = MEM[42377] + MEM[42479];
assign MEM[46121] = MEM[42378] + MEM[42402];
assign MEM[46122] = MEM[42380] + MEM[42506];
assign MEM[46123] = MEM[42384] + MEM[42427];
assign MEM[46124] = MEM[42388] + MEM[42487];
assign MEM[46125] = MEM[42389] + MEM[42420];
assign MEM[46126] = MEM[42390] + MEM[42530];
assign MEM[46127] = MEM[42392] + MEM[42516];
assign MEM[46128] = MEM[42394] + MEM[42444];
assign MEM[46129] = MEM[42395] + MEM[42493];
assign MEM[46130] = MEM[42397] + MEM[42459];
assign MEM[46131] = MEM[42398] + MEM[42496];
assign MEM[46132] = MEM[42399] + MEM[42476];
assign MEM[46133] = MEM[42400] + MEM[42442];
assign MEM[46134] = MEM[42401] + MEM[42502];
assign MEM[46135] = MEM[42403] + MEM[42448];
assign MEM[46136] = MEM[42406] + MEM[42468];
assign MEM[46137] = MEM[42407] + MEM[42424];
assign MEM[46138] = MEM[42410] + MEM[42540];
assign MEM[46139] = MEM[42411] + MEM[42467];
assign MEM[46140] = MEM[42413] + MEM[42511];
assign MEM[46141] = MEM[42415] + MEM[42537];
assign MEM[46142] = MEM[42416] + MEM[42452];
assign MEM[46143] = MEM[42417] + MEM[42491];
assign MEM[46144] = MEM[42422] + MEM[42441];
assign MEM[46145] = MEM[42423] + MEM[42503];
assign MEM[46146] = MEM[42426] + MEM[42495];
assign MEM[46147] = MEM[42428] + MEM[42473];
assign MEM[46148] = MEM[42430] + MEM[42523];
assign MEM[46149] = MEM[42431] + MEM[42462];
assign MEM[46150] = MEM[42434] + MEM[42464];
assign MEM[46151] = MEM[42435] + MEM[42509];
assign MEM[46152] = MEM[42436] + MEM[42498];
assign MEM[46153] = MEM[42438] + MEM[42472];
assign MEM[46154] = MEM[42439] + MEM[42465];
assign MEM[46155] = MEM[42440] + MEM[42541];
assign MEM[46156] = MEM[42443] + MEM[42507];
assign MEM[46157] = MEM[42446] + MEM[42510];
assign MEM[46158] = MEM[42447] + MEM[42488];
assign MEM[46159] = MEM[42449] + MEM[42527];
assign MEM[46160] = MEM[42450] + MEM[42517];
assign MEM[46161] = MEM[42451] + MEM[42549];
assign MEM[46162] = MEM[42453] + MEM[42484];
assign MEM[46163] = MEM[42455] + MEM[42463];
assign MEM[46164] = MEM[42456] + MEM[42567];
assign MEM[46165] = MEM[42457] + MEM[42481];
assign MEM[46166] = MEM[42458] + MEM[42522];
assign MEM[46167] = MEM[42461] + MEM[42535];
assign MEM[46168] = MEM[42466] + MEM[42490];
assign MEM[46169] = MEM[42470] + MEM[42550];
assign MEM[46170] = MEM[42471] + MEM[42553];
assign MEM[46171] = MEM[42474] + MEM[42500];
assign MEM[46172] = MEM[42475] + MEM[42536];
assign MEM[46173] = MEM[42477] + MEM[42560];
assign MEM[46174] = MEM[42478] + MEM[42501];
assign MEM[46175] = MEM[42480] + MEM[42532];
assign MEM[46176] = MEM[42482] + MEM[42514];
assign MEM[46177] = MEM[42483] + MEM[42561];
assign MEM[46178] = MEM[42485] + MEM[42545];
assign MEM[46179] = MEM[42486] + MEM[42534];
assign MEM[46180] = MEM[42489] + MEM[42519];
assign MEM[46181] = MEM[42492] + MEM[42539];
assign MEM[46182] = MEM[42494] + MEM[42554];
assign MEM[46183] = MEM[42497] + MEM[42607];
assign MEM[46184] = MEM[42499] + MEM[42555];
assign MEM[46185] = MEM[42504] + MEM[42508];
assign MEM[46186] = MEM[42505] + MEM[42551];
assign MEM[46187] = MEM[42512] + MEM[42574];
assign MEM[46188] = MEM[42513] + MEM[42604];
assign MEM[46189] = MEM[42515] + MEM[42562];
assign MEM[46190] = MEM[42518] + MEM[42572];
assign MEM[46191] = MEM[42520] + MEM[42584];
assign MEM[46192] = MEM[42521] + MEM[42573];
assign MEM[46193] = MEM[42524] + MEM[42615];
assign MEM[46194] = MEM[42525] + MEM[42578];
assign MEM[46195] = MEM[42526] + MEM[42595];
assign MEM[46196] = MEM[42528] + MEM[42613];
assign MEM[46197] = MEM[42529] + MEM[42602];
assign MEM[46198] = MEM[42531] + MEM[42641];
assign MEM[46199] = MEM[42533] + MEM[42565];
assign MEM[46200] = MEM[42538] + MEM[42587];
assign MEM[46201] = MEM[42542] + MEM[42556];
assign MEM[46202] = MEM[42543] + MEM[42569];
assign MEM[46203] = MEM[42544] + MEM[42601];
assign MEM[46204] = MEM[42546] + MEM[42593];
assign MEM[46205] = MEM[42547] + MEM[42617];
assign MEM[46206] = MEM[42548] + MEM[42657];
assign MEM[46207] = MEM[42552] + MEM[42616];
assign MEM[46208] = MEM[42557] + MEM[42609];
assign MEM[46209] = MEM[42558] + MEM[42681];
assign MEM[46210] = MEM[42559] + MEM[42650];
assign MEM[46211] = MEM[42563] + MEM[42605];
assign MEM[46212] = MEM[42564] + MEM[42590];
assign MEM[46213] = MEM[42566] + MEM[42610];
assign MEM[46214] = MEM[42568] + MEM[42695];
assign MEM[46215] = MEM[42570] + MEM[42647];
assign MEM[46216] = MEM[42571] + MEM[42655];
assign MEM[46217] = MEM[42575] + MEM[42634];
assign MEM[46218] = MEM[42576] + MEM[42611];
assign MEM[46219] = MEM[42577] + MEM[42589];
assign MEM[46220] = MEM[42579] + MEM[42618];
assign MEM[46221] = MEM[42580] + MEM[42598];
assign MEM[46222] = MEM[42581] + MEM[42652];
assign MEM[46223] = MEM[42582] + MEM[42637];
assign MEM[46224] = MEM[42583] + MEM[42703];
assign MEM[46225] = MEM[42585] + MEM[42643];
assign MEM[46226] = MEM[42586] + MEM[42645];
assign MEM[46227] = MEM[42588] + MEM[42674];
assign MEM[46228] = MEM[42591] + MEM[42669];
assign MEM[46229] = MEM[42592] + MEM[42659];
assign MEM[46230] = MEM[42594] + MEM[42642];
assign MEM[46231] = MEM[42596] + MEM[42718];
assign MEM[46232] = MEM[42597] + MEM[42646];
assign MEM[46233] = MEM[42599] + MEM[42683];
assign MEM[46234] = MEM[42600] + MEM[42653];
assign MEM[46235] = MEM[42603] + MEM[42640];
assign MEM[46236] = MEM[42606] + MEM[42701];
assign MEM[46237] = MEM[42608] + MEM[42633];
assign MEM[46238] = MEM[42612] + MEM[42689];
assign MEM[46239] = MEM[42614] + MEM[42742];
assign MEM[46240] = MEM[42619] + MEM[42690];
assign MEM[46241] = MEM[42620] + MEM[42687];
assign MEM[46242] = MEM[42621] + MEM[42698];
assign MEM[46243] = MEM[42622] + MEM[42716];
assign MEM[46244] = MEM[42623] + MEM[42694];
assign MEM[46245] = MEM[42624] + MEM[42649];
assign MEM[46246] = MEM[42625] + MEM[42679];
assign MEM[46247] = MEM[42626] + MEM[42665];
assign MEM[46248] = MEM[42627] + MEM[42702];
assign MEM[46249] = MEM[42628] + MEM[42715];
assign MEM[46250] = MEM[42629] + MEM[42668];
assign MEM[46251] = MEM[42630] + MEM[42661];
assign MEM[46252] = MEM[42631] + MEM[42849];
assign MEM[46253] = MEM[42632] + MEM[42662];
assign MEM[46254] = MEM[42635] + MEM[42706];
assign MEM[46255] = MEM[42636] + MEM[42763];
assign MEM[46256] = MEM[42638] + MEM[42699];
assign MEM[46257] = MEM[42639] + MEM[42744];
assign MEM[46258] = MEM[42644] + MEM[42697];
assign MEM[46259] = MEM[42648] + MEM[42712];
assign MEM[46260] = MEM[42651] + MEM[42684];
assign MEM[46261] = MEM[42654] + MEM[42696];
assign MEM[46262] = MEM[42656] + MEM[42731];
assign MEM[46263] = MEM[42658] + MEM[42686];
assign MEM[46264] = MEM[42660] + MEM[42709];
assign MEM[46265] = MEM[42663] + MEM[42729];
assign MEM[46266] = MEM[42664] + MEM[42812];
assign MEM[46267] = MEM[42666] + MEM[42692];
assign MEM[46268] = MEM[42667] + MEM[42727];
assign MEM[46269] = MEM[42670] + MEM[42734];
assign MEM[46270] = MEM[42671] + MEM[42688];
assign MEM[46271] = MEM[42672] + MEM[42723];
assign MEM[46272] = MEM[42673] + MEM[42746];
assign MEM[46273] = MEM[42675] + MEM[42789];
assign MEM[46274] = MEM[42676] + MEM[42738];
assign MEM[46275] = MEM[42677] + MEM[42769];
assign MEM[46276] = MEM[42678] + MEM[42720];
assign MEM[46277] = MEM[42680] + MEM[42743];
assign MEM[46278] = MEM[42682] + MEM[42736];
assign MEM[46279] = MEM[42685] + MEM[42757];
assign MEM[46280] = MEM[42691] + MEM[42760];
assign MEM[46281] = MEM[42693] + MEM[42779];
assign MEM[46282] = MEM[42700] + MEM[42710];
assign MEM[46283] = MEM[42704] + MEM[42793];
assign MEM[46284] = MEM[42705] + MEM[42780];
assign MEM[46285] = MEM[42707] + MEM[42813];
assign MEM[46286] = MEM[42708] + MEM[42739];
assign MEM[46287] = MEM[42711] + MEM[42784];
assign MEM[46288] = MEM[42713] + MEM[42753];
assign MEM[46289] = MEM[42714] + MEM[42782];
assign MEM[46290] = MEM[42717] + MEM[42795];
assign MEM[46291] = MEM[42719] + MEM[42798];
assign MEM[46292] = MEM[42721] + MEM[42772];
assign MEM[46293] = MEM[42722] + MEM[42771];
assign MEM[46294] = MEM[42724] + MEM[42808];
assign MEM[46295] = MEM[42725] + MEM[42806];
assign MEM[46296] = MEM[42726] + MEM[42735];
assign MEM[46297] = MEM[42728] + MEM[42809];
assign MEM[46298] = MEM[42730] + MEM[42759];
assign MEM[46299] = MEM[42732] + MEM[42824];
assign MEM[46300] = MEM[42733] + MEM[42775];
assign MEM[46301] = MEM[42737] + MEM[42777];
assign MEM[46302] = MEM[42740] + MEM[42801];
assign MEM[46303] = MEM[42741] + MEM[42855];
assign MEM[46304] = MEM[42745] + MEM[42810];
assign MEM[46305] = MEM[42747] + MEM[42815];
assign MEM[46306] = MEM[42748] + MEM[42817];
assign MEM[46307] = MEM[42749] + MEM[42799];
assign MEM[46308] = MEM[42750] + MEM[42807];
assign MEM[46309] = MEM[42751] + MEM[42821];
assign MEM[46310] = MEM[42752] + MEM[42791];
assign MEM[46311] = MEM[42754] + MEM[42773];
assign MEM[46312] = MEM[42755] + MEM[42786];
assign MEM[46313] = MEM[42756] + MEM[42835];
assign MEM[46314] = MEM[42758] + MEM[42814];
assign MEM[46315] = MEM[42761] + MEM[42820];
assign MEM[46316] = MEM[42762] + MEM[42800];
assign MEM[46317] = MEM[42764] + MEM[42929];
assign MEM[46318] = MEM[42765] + MEM[42941];
assign MEM[46319] = MEM[42766] + MEM[42864];
assign MEM[46320] = MEM[42767] + MEM[42896];
assign MEM[46321] = MEM[42768] + MEM[42826];
assign MEM[46322] = MEM[42770] + MEM[42805];
assign MEM[46323] = MEM[42774] + MEM[42840];
assign MEM[46324] = MEM[42776] + MEM[42832];
assign MEM[46325] = MEM[42778] + MEM[42869];
assign MEM[46326] = MEM[42781] + MEM[42839];
assign MEM[46327] = MEM[42783] + MEM[42827];
assign MEM[46328] = MEM[42785] + MEM[42833];
assign MEM[46329] = MEM[42787] + MEM[42825];
assign MEM[46330] = MEM[42788] + MEM[42846];
assign MEM[46331] = MEM[42790] + MEM[42856];
assign MEM[46332] = MEM[42792] + MEM[42949];
assign MEM[46333] = MEM[42794] + MEM[42830];
assign MEM[46334] = MEM[42796] + MEM[42816];
assign MEM[46335] = MEM[42797] + MEM[42853];
assign MEM[46336] = MEM[42802] + MEM[42837];
assign MEM[46337] = MEM[42803] + MEM[42822];
assign MEM[46338] = MEM[42804] + MEM[42851];
assign MEM[46339] = MEM[42811] + MEM[42894];
assign MEM[46340] = MEM[42818] + MEM[42841];
assign MEM[46341] = MEM[42819] + MEM[42854];
assign MEM[46342] = MEM[42823] + MEM[42865];
assign MEM[46343] = MEM[42828] + MEM[42883];
assign MEM[46344] = MEM[42829] + MEM[42915];
assign MEM[46345] = MEM[42831] + MEM[42863];
assign MEM[46346] = MEM[42834] + MEM[42892];
assign MEM[46347] = MEM[42836] + MEM[42990];
assign MEM[46348] = MEM[42838] + MEM[42875];
assign MEM[46349] = MEM[42842] + MEM[42928];
assign MEM[46350] = MEM[42843] + MEM[42913];
assign MEM[46351] = MEM[42844] + MEM[42919];
assign MEM[46352] = MEM[42845] + MEM[42910];
assign MEM[46353] = MEM[42847] + MEM[42901];
assign MEM[46354] = MEM[42848] + MEM[42918];
assign MEM[46355] = MEM[42850] + MEM[42870];
assign MEM[46356] = MEM[42852] + MEM[42882];
assign MEM[46357] = MEM[42857] + MEM[42925];
assign MEM[46358] = MEM[42858] + MEM[42898];
assign MEM[46359] = MEM[42859] + MEM[42886];
assign MEM[46360] = MEM[42860] + MEM[42905];
assign MEM[46361] = MEM[42861] + MEM[42924];
assign MEM[46362] = MEM[42862] + MEM[42943];
assign MEM[46363] = MEM[42866] + MEM[42931];
assign MEM[46364] = MEM[42867] + MEM[42922];
assign MEM[46365] = MEM[42868] + MEM[42917];
assign MEM[46366] = MEM[42871] + MEM[42906];
assign MEM[46367] = MEM[42872] + MEM[42936];
assign MEM[46368] = MEM[42873] + MEM[42891];
assign MEM[46369] = MEM[42874] + MEM[42967];
assign MEM[46370] = MEM[42876] + MEM[42902];
assign MEM[46371] = MEM[42877] + MEM[42908];
assign MEM[46372] = MEM[42878] + MEM[43017];
assign MEM[46373] = MEM[42879] + MEM[42947];
assign MEM[46374] = MEM[42880] + MEM[42951];
assign MEM[46375] = MEM[42881] + MEM[42997];
assign MEM[46376] = MEM[42884] + MEM[43040];
assign MEM[46377] = MEM[42885] + MEM[42933];
assign MEM[46378] = MEM[42887] + MEM[42944];
assign MEM[46379] = MEM[42888] + MEM[42969];
assign MEM[46380] = MEM[42889] + MEM[42946];
assign MEM[46381] = MEM[42890] + MEM[42993];
assign MEM[46382] = MEM[42893] + MEM[42945];
assign MEM[46383] = MEM[42895] + MEM[42955];
assign MEM[46384] = MEM[42897] + MEM[42953];
assign MEM[46385] = MEM[42899] + MEM[42940];
assign MEM[46386] = MEM[42900] + MEM[42982];
assign MEM[46387] = MEM[42903] + MEM[42952];
assign MEM[46388] = MEM[42904] + MEM[42942];
assign MEM[46389] = MEM[42907] + MEM[42978];
assign MEM[46390] = MEM[42909] + MEM[42959];
assign MEM[46391] = MEM[42911] + MEM[42939];
assign MEM[46392] = MEM[42912] + MEM[42975];
assign MEM[46393] = MEM[42914] + MEM[43004];
assign MEM[46394] = MEM[42916] + MEM[43001];
assign MEM[46395] = MEM[42920] + MEM[42994];
assign MEM[46396] = MEM[42921] + MEM[42956];
assign MEM[46397] = MEM[42923] + MEM[43015];
assign MEM[46398] = MEM[42926] + MEM[42974];
assign MEM[46399] = MEM[42927] + MEM[42957];
assign MEM[46400] = MEM[42930] + MEM[42960];
assign MEM[46401] = MEM[42932] + MEM[43039];
assign MEM[46402] = MEM[42934] + MEM[43035];
assign MEM[46403] = MEM[42935] + MEM[43012];
assign MEM[46404] = MEM[42937] + MEM[42966];
assign MEM[46405] = MEM[42938] + MEM[42977];
assign MEM[46406] = MEM[42948] + MEM[43014];
assign MEM[46407] = MEM[42950] + MEM[43026];
assign MEM[46408] = MEM[42954] + MEM[42991];
assign MEM[46409] = MEM[42958] + MEM[42989];
assign MEM[46410] = MEM[42961] + MEM[43034];
assign MEM[46411] = MEM[42962] + MEM[43013];
assign MEM[46412] = MEM[42963] + MEM[43073];
assign MEM[46413] = MEM[42964] + MEM[42985];
assign MEM[46414] = MEM[42965] + MEM[42987];
assign MEM[46415] = MEM[42968] + MEM[43025];
assign MEM[46416] = MEM[42970] + MEM[43067];
assign MEM[46417] = MEM[42971] + MEM[43045];
assign MEM[46418] = MEM[42972] + MEM[43010];
assign MEM[46419] = MEM[42973] + MEM[43047];
assign MEM[46420] = MEM[42976] + MEM[43016];
assign MEM[46421] = MEM[42979] + MEM[43058];
assign MEM[46422] = MEM[42980] + MEM[43108];
assign MEM[46423] = MEM[42981] + MEM[43057];
assign MEM[46424] = MEM[42983] + MEM[43022];
assign MEM[46425] = MEM[42984] + MEM[43018];
assign MEM[46426] = MEM[42986] + MEM[43038];
assign MEM[46427] = MEM[42988] + MEM[43020];
assign MEM[46428] = MEM[42992] + MEM[43068];
assign MEM[46429] = MEM[42995] + MEM[43093];
assign MEM[46430] = MEM[42996] + MEM[43097];
assign MEM[46431] = MEM[42998] + MEM[43048];
assign MEM[46432] = MEM[42999] + MEM[43055];
assign MEM[46433] = MEM[43000] + MEM[43066];
assign MEM[46434] = MEM[43002] + MEM[43029];
assign MEM[46435] = MEM[43003] + MEM[43062];
assign MEM[46436] = MEM[43005] + MEM[43098];
assign MEM[46437] = MEM[43006] + MEM[43028];
assign MEM[46438] = MEM[43007] + MEM[43051];
assign MEM[46439] = MEM[43008] + MEM[43076];
assign MEM[46440] = MEM[43009] + MEM[43046];
assign MEM[46441] = MEM[43011] + MEM[43085];
assign MEM[46442] = MEM[43019] + MEM[43117];
assign MEM[46443] = MEM[43021] + MEM[43078];
assign MEM[46444] = MEM[43023] + MEM[43074];
assign MEM[46445] = MEM[43024] + MEM[43081];
assign MEM[46446] = MEM[43027] + MEM[43052];
assign MEM[46447] = MEM[43030] + MEM[43114];
assign MEM[46448] = MEM[43031] + MEM[43091];
assign MEM[46449] = MEM[43032] + MEM[43087];
assign MEM[46450] = MEM[43033] + MEM[43111];
assign MEM[46451] = MEM[43036] + MEM[43104];
assign MEM[46452] = MEM[43037] + MEM[43126];
assign MEM[46453] = MEM[43041] + MEM[43089];
assign MEM[46454] = MEM[43042] + MEM[43103];
assign MEM[46455] = MEM[43043] + MEM[43065];
assign MEM[46456] = MEM[43044] + MEM[43116];
assign MEM[46457] = MEM[43049] + MEM[43124];
assign MEM[46458] = MEM[43050] + MEM[43086];
assign MEM[46459] = MEM[43053] + MEM[43082];
assign MEM[46460] = MEM[43054] + MEM[43105];
assign MEM[46461] = MEM[43056] + MEM[43145];
assign MEM[46462] = MEM[43059] + MEM[43118];
assign MEM[46463] = MEM[43060] + MEM[43110];
assign MEM[46464] = MEM[43061] + MEM[43123];
assign MEM[46465] = MEM[43063] + MEM[43142];
assign MEM[46466] = MEM[43064] + MEM[43119];
assign MEM[46467] = MEM[43069] + MEM[43138];
assign MEM[46468] = MEM[43070] + MEM[43080];
assign MEM[46469] = MEM[43071] + MEM[43112];
assign MEM[46470] = MEM[43072] + MEM[43096];
assign MEM[46471] = MEM[43075] + MEM[43162];
assign MEM[46472] = MEM[43077] + MEM[43115];
assign MEM[46473] = MEM[43079] + MEM[43171];
assign MEM[46474] = MEM[43083] + MEM[43127];
assign MEM[46475] = MEM[43084] + MEM[43158];
assign MEM[46476] = MEM[43088] + MEM[43189];
assign MEM[46477] = MEM[43090] + MEM[43267];
assign MEM[46478] = MEM[43092] + MEM[43209];
assign MEM[46479] = MEM[43094] + MEM[43191];
assign MEM[46480] = MEM[43095] + MEM[43181];
assign MEM[46481] = MEM[43099] + MEM[43168];
assign MEM[46482] = MEM[43100] + MEM[43212];
assign MEM[46483] = MEM[43101] + MEM[43182];
assign MEM[46484] = MEM[43102] + MEM[43166];
assign MEM[46485] = MEM[43106] + MEM[43150];
assign MEM[46486] = MEM[43107] + MEM[43232];
assign MEM[46487] = MEM[43109] + MEM[43202];
assign MEM[46488] = MEM[43113] + MEM[43190];
assign MEM[46489] = MEM[43120] + MEM[43155];
assign MEM[46490] = MEM[43121] + MEM[43161];
assign MEM[46491] = MEM[43122] + MEM[43169];
assign MEM[46492] = MEM[43125] + MEM[43157];
assign MEM[46493] = MEM[43128] + MEM[43203];
assign MEM[46494] = MEM[43129] + MEM[43167];
assign MEM[46495] = MEM[43130] + MEM[43215];
assign MEM[46496] = MEM[43131] + MEM[43177];
assign MEM[46497] = MEM[43132] + MEM[43176];
assign MEM[46498] = MEM[43133] + MEM[43338];
assign MEM[46499] = MEM[43134] + MEM[43205];
assign MEM[46500] = MEM[43135] + MEM[43260];
assign MEM[46501] = MEM[43136] + MEM[43239];
assign MEM[46502] = MEM[43137] + MEM[43235];
assign MEM[46503] = MEM[43139] + MEM[43185];
assign MEM[46504] = MEM[43140] + MEM[43247];
assign MEM[46505] = MEM[43141] + MEM[43201];
assign MEM[46506] = MEM[43143] + MEM[43187];
assign MEM[46507] = MEM[43144] + MEM[43204];
assign MEM[46508] = MEM[43146] + MEM[43246];
assign MEM[46509] = MEM[43147] + MEM[43225];
assign MEM[46510] = MEM[43148] + MEM[43188];
assign MEM[46511] = MEM[43149] + MEM[43173];
assign MEM[46512] = MEM[43151] + MEM[43217];
assign MEM[46513] = MEM[43152] + MEM[43206];
assign MEM[46514] = MEM[43153] + MEM[43178];
assign MEM[46515] = MEM[43154] + MEM[43224];
assign MEM[46516] = MEM[43156] + MEM[43227];
assign MEM[46517] = MEM[43159] + MEM[43323];
assign MEM[46518] = MEM[43160] + MEM[43251];
assign MEM[46519] = MEM[43163] + MEM[43277];
assign MEM[46520] = MEM[43164] + MEM[43253];
assign MEM[46521] = MEM[43165] + MEM[43244];
assign MEM[46522] = MEM[43170] + MEM[43219];
assign MEM[46523] = MEM[43172] + MEM[43194];
assign MEM[46524] = MEM[43174] + MEM[43252];
assign MEM[46525] = MEM[43175] + MEM[43210];
assign MEM[46526] = MEM[43179] + MEM[43193];
assign MEM[46527] = MEM[43180] + MEM[43339];
assign MEM[46528] = MEM[43183] + MEM[43234];
assign MEM[46529] = MEM[43184] + MEM[43294];
assign MEM[46530] = MEM[43186] + MEM[43236];
assign MEM[46531] = MEM[43192] + MEM[43375];
assign MEM[46532] = MEM[43195] + MEM[43271];
assign MEM[46533] = MEM[43196] + MEM[43222];
assign MEM[46534] = MEM[43197] + MEM[43318];
assign MEM[46535] = MEM[43198] + MEM[43283];
assign MEM[46536] = MEM[43199] + MEM[43254];
assign MEM[46537] = MEM[43200] + MEM[43218];
assign MEM[46538] = MEM[43207] + MEM[43296];
assign MEM[46539] = MEM[43208] + MEM[43276];
assign MEM[46540] = MEM[43211] + MEM[43242];
assign MEM[46541] = MEM[43213] + MEM[43257];
assign MEM[46542] = MEM[43214] + MEM[43303];
assign MEM[46543] = MEM[43216] + MEM[43249];
assign MEM[46544] = MEM[43220] + MEM[43273];
assign MEM[46545] = MEM[43221] + MEM[43295];
assign MEM[46546] = MEM[43223] + MEM[43269];
assign MEM[46547] = MEM[43226] + MEM[43301];
assign MEM[46548] = MEM[43228] + MEM[43386];
assign MEM[46549] = MEM[43229] + MEM[43248];
assign MEM[46550] = MEM[43230] + MEM[43261];
assign MEM[46551] = MEM[43231] + MEM[43266];
assign MEM[46552] = MEM[43233] + MEM[43321];
assign MEM[46553] = MEM[43237] + MEM[43354];
assign MEM[46554] = MEM[43238] + MEM[43286];
assign MEM[46555] = MEM[43240] + MEM[43280];
assign MEM[46556] = MEM[43241] + MEM[43290];
assign MEM[46557] = MEM[43243] + MEM[43278];
assign MEM[46558] = MEM[43245] + MEM[43291];
assign MEM[46559] = MEM[43250] + MEM[43311];
assign MEM[46560] = MEM[43255] + MEM[43324];
assign MEM[46561] = MEM[43256] + MEM[43305];
assign MEM[46562] = MEM[43258] + MEM[43293];
assign MEM[46563] = MEM[43259] + MEM[43334];
assign MEM[46564] = MEM[43262] + MEM[43345];
assign MEM[46565] = MEM[43263] + MEM[43418];
assign MEM[46566] = MEM[43264] + MEM[43320];
assign MEM[46567] = MEM[43265] + MEM[43299];
assign MEM[46568] = MEM[43268] + MEM[43355];
assign MEM[46569] = MEM[43270] + MEM[43333];
assign MEM[46570] = MEM[43272] + MEM[43298];
assign MEM[46571] = MEM[43274] + MEM[43325];
assign MEM[46572] = MEM[43275] + MEM[43317];
assign MEM[46573] = MEM[43279] + MEM[43332];
assign MEM[46574] = MEM[43281] + MEM[43330];
assign MEM[46575] = MEM[43282] + MEM[43357];
assign MEM[46576] = MEM[43284] + MEM[43346];
assign MEM[46577] = MEM[43285] + MEM[43316];
assign MEM[46578] = MEM[43287] + MEM[43358];
assign MEM[46579] = MEM[43288] + MEM[43382];
assign MEM[46580] = MEM[43289] + MEM[43363];
assign MEM[46581] = MEM[43292] + MEM[43319];
assign MEM[46582] = MEM[43297] + MEM[43348];
assign MEM[46583] = MEM[43300] + MEM[43350];
assign MEM[46584] = MEM[43302] + MEM[43380];
assign MEM[46585] = MEM[43304] + MEM[43351];
assign MEM[46586] = MEM[43306] + MEM[43360];
assign MEM[46587] = MEM[43307] + MEM[43361];
assign MEM[46588] = MEM[43308] + MEM[43322];
assign MEM[46589] = MEM[43309] + MEM[43344];
assign MEM[46590] = MEM[43310] + MEM[43384];
assign MEM[46591] = MEM[43312] + MEM[43393];
assign MEM[46592] = MEM[43313] + MEM[43368];
assign MEM[46593] = MEM[43314] + MEM[43397];
assign MEM[46594] = MEM[43315] + MEM[43366];
assign MEM[46595] = MEM[43326] + MEM[43369];
assign MEM[46596] = MEM[43327] + MEM[43367];
assign MEM[46597] = MEM[43328] + MEM[43335];
assign MEM[46598] = MEM[43329] + MEM[43388];
assign MEM[46599] = MEM[43331] + MEM[43432];
assign MEM[46600] = MEM[43336] + MEM[43429];
assign MEM[46601] = MEM[43337] + MEM[43434];
assign MEM[46602] = MEM[43340] + MEM[43456];
assign MEM[46603] = MEM[43341] + MEM[43454];
assign MEM[46604] = MEM[43342] + MEM[43401];
assign MEM[46605] = MEM[43343] + MEM[43395];
assign MEM[46606] = MEM[43347] + MEM[43464];
assign MEM[46607] = MEM[43349] + MEM[43376];
assign MEM[46608] = MEM[43352] + MEM[43427];
assign MEM[46609] = MEM[43353] + MEM[43412];
assign MEM[46610] = MEM[43356] + MEM[43373];
assign MEM[46611] = MEM[43359] + MEM[43371];
assign MEM[46612] = MEM[43362] + MEM[43446];
assign MEM[46613] = MEM[43364] + MEM[43392];
assign MEM[46614] = MEM[43365] + MEM[43414];
assign MEM[46615] = MEM[43370] + MEM[43396];
assign MEM[46616] = MEM[43372] + MEM[43428];
assign MEM[46617] = MEM[43374] + MEM[43453];
assign MEM[46618] = MEM[43377] + MEM[43424];
assign MEM[46619] = MEM[43378] + MEM[43440];
assign MEM[46620] = MEM[43379] + MEM[43436];
assign MEM[46621] = MEM[43381] + MEM[43496];
assign MEM[46622] = MEM[43383] + MEM[43462];
assign MEM[46623] = MEM[43385] + MEM[43473];
assign MEM[46624] = MEM[43387] + MEM[43495];
assign MEM[46625] = MEM[43389] + MEM[43422];
assign MEM[46626] = MEM[43390] + MEM[43439];
assign MEM[46627] = MEM[43391] + MEM[43490];
assign MEM[46628] = MEM[43394] + MEM[43444];
assign MEM[46629] = MEM[43398] + MEM[43524];
assign MEM[46630] = MEM[43399] + MEM[43475];
assign MEM[46631] = MEM[43400] + MEM[43511];
assign MEM[46632] = MEM[43402] + MEM[43435];
assign MEM[46633] = MEM[43403] + MEM[43478];
assign MEM[46634] = MEM[43404] + MEM[43433];
assign MEM[46635] = MEM[43405] + MEM[43455];
assign MEM[46636] = MEM[43406] + MEM[43447];
assign MEM[46637] = MEM[43407] + MEM[43460];
assign MEM[46638] = MEM[43408] + MEM[43437];
assign MEM[46639] = MEM[43409] + MEM[43501];
assign MEM[46640] = MEM[43410] + MEM[43505];
assign MEM[46641] = MEM[43411] + MEM[43477];
assign MEM[46642] = MEM[43413] + MEM[43470];
assign MEM[46643] = MEM[43415] + MEM[43479];
assign MEM[46644] = MEM[43416] + MEM[43543];
assign MEM[46645] = MEM[43417] + MEM[43474];
assign MEM[46646] = MEM[43419] + MEM[43482];
assign MEM[46647] = MEM[43420] + MEM[43451];
assign MEM[46648] = MEM[43421] + MEM[43510];
assign MEM[46649] = MEM[43423] + MEM[43558];
assign MEM[46650] = MEM[43425] + MEM[43507];
assign MEM[46651] = MEM[43426] + MEM[43522];
assign MEM[46652] = MEM[43430] + MEM[43489];
assign MEM[46653] = MEM[43431] + MEM[43461];
assign MEM[46654] = MEM[43438] + MEM[43463];
assign MEM[46655] = MEM[43441] + MEM[43497];
assign MEM[46656] = MEM[43442] + MEM[43518];
assign MEM[46657] = MEM[43443] + MEM[43551];
assign MEM[46658] = MEM[43445] + MEM[43506];
assign MEM[46659] = MEM[43448] + MEM[43540];
assign MEM[46660] = MEM[43449] + MEM[43537];
assign MEM[46661] = MEM[43450] + MEM[43559];
assign MEM[46662] = MEM[43452] + MEM[43466];
assign MEM[46663] = MEM[43457] + MEM[43500];
assign MEM[46664] = MEM[43458] + MEM[43498];
assign MEM[46665] = MEM[43459] + MEM[43488];
assign MEM[46666] = MEM[43465] + MEM[43572];
assign MEM[46667] = MEM[43467] + MEM[43556];
assign MEM[46668] = MEM[43468] + MEM[43548];
assign MEM[46669] = MEM[43469] + MEM[43514];
assign MEM[46670] = MEM[43471] + MEM[43571];
assign MEM[46671] = MEM[43472] + MEM[43492];
assign MEM[46672] = MEM[43476] + MEM[43520];
assign MEM[46673] = MEM[43480] + MEM[43502];
assign MEM[46674] = MEM[43481] + MEM[43487];
assign MEM[46675] = MEM[43483] + MEM[43557];
assign MEM[46676] = MEM[43484] + MEM[43538];
assign MEM[46677] = MEM[43485] + MEM[43513];
assign MEM[46678] = MEM[43486] + MEM[43561];
assign MEM[46679] = MEM[43491] + MEM[43570];
assign MEM[46680] = MEM[43493] + MEM[43544];
assign MEM[46681] = MEM[43494] + MEM[43516];
assign MEM[46682] = MEM[43499] + MEM[43575];
assign MEM[46683] = MEM[43503] + MEM[43547];
assign MEM[46684] = MEM[43504] + MEM[43532];
assign MEM[46685] = MEM[43508] + MEM[43582];
assign MEM[46686] = MEM[43509] + MEM[43603];
assign MEM[46687] = MEM[43512] + MEM[43567];
assign MEM[46688] = MEM[43515] + MEM[43560];
assign MEM[46689] = MEM[43517] + MEM[43529];
assign MEM[46690] = MEM[43519] + MEM[43552];
assign MEM[46691] = MEM[43521] + MEM[43597];
assign MEM[46692] = MEM[43523] + MEM[43638];
assign MEM[46693] = MEM[43525] + MEM[43595];
assign MEM[46694] = MEM[43526] + MEM[43607];
assign MEM[46695] = MEM[43527] + MEM[43565];
assign MEM[46696] = MEM[43528] + MEM[43586];
assign MEM[46697] = MEM[43530] + MEM[43568];
assign MEM[46698] = MEM[43531] + MEM[43609];
assign MEM[46699] = MEM[43533] + MEM[43605];
assign MEM[46700] = MEM[43534] + MEM[43574];
assign MEM[46701] = MEM[43535] + MEM[43576];
assign MEM[46702] = MEM[43536] + MEM[43720];
assign MEM[46703] = MEM[43539] + MEM[43602];
assign MEM[46704] = MEM[43541] + MEM[43606];
assign MEM[46705] = MEM[43542] + MEM[43584];
assign MEM[46706] = MEM[43545] + MEM[43685];
assign MEM[46707] = MEM[43546] + MEM[43578];
assign MEM[46708] = MEM[43549] + MEM[43573];
assign MEM[46709] = MEM[43550] + MEM[43663];
assign MEM[46710] = MEM[43553] + MEM[43580];
assign MEM[46711] = MEM[43554] + MEM[43634];
assign MEM[46712] = MEM[43555] + MEM[43683];
assign MEM[46713] = MEM[43562] + MEM[43598];
assign MEM[46714] = MEM[43563] + MEM[43635];
assign MEM[46715] = MEM[43564] + MEM[43664];
assign MEM[46716] = MEM[43566] + MEM[43594];
assign MEM[46717] = MEM[43569] + MEM[43633];
assign MEM[46718] = MEM[43577] + MEM[43630];
assign MEM[46719] = MEM[43579] + MEM[43614];
assign MEM[46720] = MEM[43581] + MEM[43610];
assign MEM[46721] = MEM[43583] + MEM[43655];
assign MEM[46722] = MEM[43585] + MEM[43719];
assign MEM[46723] = MEM[43587] + MEM[43665];
assign MEM[46724] = MEM[43588] + MEM[43680];
assign MEM[46725] = MEM[43589] + MEM[43707];
assign MEM[46726] = MEM[43590] + MEM[43617];
assign MEM[46727] = MEM[43591] + MEM[43651];
assign MEM[46728] = MEM[43592] + MEM[43670];
assign MEM[46729] = MEM[43593] + MEM[43672];
assign MEM[46730] = MEM[43596] + MEM[43637];
assign MEM[46731] = MEM[43599] + MEM[43640];
assign MEM[46732] = MEM[43600] + MEM[43699];
assign MEM[46733] = MEM[43601] + MEM[43682];
assign MEM[46734] = MEM[43604] + MEM[43717];
assign MEM[46735] = MEM[43608] + MEM[43652];
assign MEM[46736] = MEM[43611] + MEM[43628];
assign MEM[46737] = MEM[43612] + MEM[43632];
assign MEM[46738] = MEM[43613] + MEM[43662];
assign MEM[46739] = MEM[43615] + MEM[43686];
assign MEM[46740] = MEM[43616] + MEM[43649];
assign MEM[46741] = MEM[43618] + MEM[43647];
assign MEM[46742] = MEM[43619] + MEM[43669];
assign MEM[46743] = MEM[43620] + MEM[43715];
assign MEM[46744] = MEM[43621] + MEM[43650];
assign MEM[46745] = MEM[43622] + MEM[43688];
assign MEM[46746] = MEM[43623] + MEM[43676];
assign MEM[46747] = MEM[43624] + MEM[43660];
assign MEM[46748] = MEM[43625] + MEM[43675];
assign MEM[46749] = MEM[43626] + MEM[43677];
assign MEM[46750] = MEM[43627] + MEM[43661];
assign MEM[46751] = MEM[43629] + MEM[43667];
assign MEM[46752] = MEM[43631] + MEM[43646];
assign MEM[46753] = MEM[43636] + MEM[43739];
assign MEM[46754] = MEM[43639] + MEM[43695];
assign MEM[46755] = MEM[43641] + MEM[43671];
assign MEM[46756] = MEM[43642] + MEM[43734];
assign MEM[46757] = MEM[43643] + MEM[43764];
assign MEM[46758] = MEM[43644] + MEM[43687];
assign MEM[46759] = MEM[43645] + MEM[43714];
assign MEM[46760] = MEM[43648] + MEM[43691];
assign MEM[46761] = MEM[43653] + MEM[43728];
assign MEM[46762] = MEM[43654] + MEM[43726];
assign MEM[46763] = MEM[43656] + MEM[43742];
assign MEM[46764] = MEM[43657] + MEM[43703];
assign MEM[46765] = MEM[43658] + MEM[43701];
assign MEM[46766] = MEM[43659] + MEM[43730];
assign MEM[46767] = MEM[43666] + MEM[43732];
assign MEM[46768] = MEM[43668] + MEM[43694];
assign MEM[46769] = MEM[43673] + MEM[43704];
assign MEM[46770] = MEM[43674] + MEM[43713];
assign MEM[46771] = MEM[43678] + MEM[43729];
assign MEM[46772] = MEM[43679] + MEM[43712];
assign MEM[46773] = MEM[43681] + MEM[43741];
assign MEM[46774] = MEM[43684] + MEM[43702];
assign MEM[46775] = MEM[43689] + MEM[43727];
assign MEM[46776] = MEM[43690] + MEM[43752];
assign MEM[46777] = MEM[43692] + MEM[43836];
assign MEM[46778] = MEM[43693] + MEM[43755];
assign MEM[46779] = MEM[43696] + MEM[43723];
assign MEM[46780] = MEM[43697] + MEM[43818];
assign MEM[46781] = MEM[43698] + MEM[43740];
assign MEM[46782] = MEM[43700] + MEM[43769];
assign MEM[46783] = MEM[43705] + MEM[43758];
assign MEM[46784] = MEM[43706] + MEM[43735];
assign MEM[46785] = MEM[43708] + MEM[43791];
assign MEM[46786] = MEM[43709] + MEM[43809];
assign MEM[46787] = MEM[43710] + MEM[43744];
assign MEM[46788] = MEM[43711] + MEM[43775];
assign MEM[46789] = MEM[43716] + MEM[43759];
assign MEM[46790] = MEM[43718] + MEM[43872];
assign MEM[46791] = MEM[43721] + MEM[43776];
assign MEM[46792] = MEM[43722] + MEM[43820];
assign MEM[46793] = MEM[43724] + MEM[43748];
assign MEM[46794] = MEM[43725] + MEM[43795];
assign MEM[46795] = MEM[43731] + MEM[43788];
assign MEM[46796] = MEM[43733] + MEM[43787];
assign MEM[46797] = MEM[43736] + MEM[43941];
assign MEM[46798] = MEM[43737] + MEM[43838];
assign MEM[46799] = MEM[43738] + MEM[43785];
assign MEM[46800] = MEM[43743] + MEM[43790];
assign MEM[46801] = MEM[43745] + MEM[43805];
assign MEM[46802] = MEM[43746] + MEM[43830];
assign MEM[46803] = MEM[43747] + MEM[43798];
assign MEM[46804] = MEM[43749] + MEM[43770];
assign MEM[46805] = MEM[43750] + MEM[43871];
assign MEM[46806] = MEM[43751] + MEM[43793];
assign MEM[46807] = MEM[43753] + MEM[43783];
assign MEM[46808] = MEM[43754] + MEM[43814];
assign MEM[46809] = MEM[43756] + MEM[43773];
assign MEM[46810] = MEM[43757] + MEM[43833];
assign MEM[46811] = MEM[43760] + MEM[43781];
assign MEM[46812] = MEM[43761] + MEM[43799];
assign MEM[46813] = MEM[43762] + MEM[43856];
assign MEM[46814] = MEM[43763] + MEM[43848];
assign MEM[46815] = MEM[43765] + MEM[43859];
assign MEM[46816] = MEM[43766] + MEM[43801];
assign MEM[46817] = MEM[43767] + MEM[43792];
assign MEM[46818] = MEM[43768] + MEM[43870];
assign MEM[46819] = MEM[43771] + MEM[43832];
assign MEM[46820] = MEM[43772] + MEM[43831];
assign MEM[46821] = MEM[43774] + MEM[43862];
assign MEM[46822] = MEM[43777] + MEM[43840];
assign MEM[46823] = MEM[43778] + MEM[43803];
assign MEM[46824] = MEM[43779] + MEM[43825];
assign MEM[46825] = MEM[43780] + MEM[43829];
assign MEM[46826] = MEM[43782] + MEM[43929];
assign MEM[46827] = MEM[43784] + MEM[43821];
assign MEM[46828] = MEM[43786] + MEM[43842];
assign MEM[46829] = MEM[43789] + MEM[43828];
assign MEM[46830] = MEM[43794] + MEM[43868];
assign MEM[46831] = MEM[43796] + MEM[43824];
assign MEM[46832] = MEM[43797] + MEM[43855];
assign MEM[46833] = MEM[43800] + MEM[43863];
assign MEM[46834] = MEM[43802] + MEM[43822];
assign MEM[46835] = MEM[43804] + MEM[43851];
assign MEM[46836] = MEM[43806] + MEM[43876];
assign MEM[46837] = MEM[43807] + MEM[43844];
assign MEM[46838] = MEM[43808] + MEM[43847];
assign MEM[46839] = MEM[43810] + MEM[43917];
assign MEM[46840] = MEM[43811] + MEM[43873];
assign MEM[46841] = MEM[43812] + MEM[43869];
assign MEM[46842] = MEM[43813] + MEM[43858];
assign MEM[46843] = MEM[43815] + MEM[43911];
assign MEM[46844] = MEM[43816] + MEM[43912];
assign MEM[46845] = MEM[43817] + MEM[43895];
assign MEM[46846] = MEM[43819] + MEM[43865];
assign MEM[46847] = MEM[43823] + MEM[43913];
assign MEM[46848] = MEM[43826] + MEM[43901];
assign MEM[46849] = MEM[43827] + MEM[43922];
assign MEM[46850] = MEM[43834] + MEM[43877];
assign MEM[46851] = MEM[43835] + MEM[43867];
assign MEM[46852] = MEM[43837] + MEM[43915];
assign MEM[46853] = MEM[43839] + MEM[43906];
assign MEM[46854] = MEM[43841] + MEM[43920];
assign MEM[46855] = MEM[43843] + MEM[43956];
assign MEM[46856] = MEM[43845] + MEM[43953];
assign MEM[46857] = MEM[43846] + MEM[43899];
assign MEM[46858] = MEM[43849] + MEM[43925];
assign MEM[46859] = MEM[43850] + MEM[43898];
assign MEM[46860] = MEM[43852] + MEM[43921];
assign MEM[46861] = MEM[43853] + MEM[43914];
assign MEM[46862] = MEM[43854] + MEM[43884];
assign MEM[46863] = MEM[43857] + MEM[43893];
assign MEM[46864] = MEM[43860] + MEM[43894];
assign MEM[46865] = MEM[43861] + MEM[43970];
assign MEM[46866] = MEM[43864] + MEM[43900];
assign MEM[46867] = MEM[43866] + MEM[43942];
assign MEM[46868] = MEM[43874] + MEM[43987];
assign MEM[46869] = MEM[43875] + MEM[43927];
assign MEM[46870] = MEM[43878] + MEM[43950];
assign MEM[46871] = MEM[43879] + MEM[43919];
assign MEM[46872] = MEM[43880] + MEM[43897];
assign MEM[46873] = MEM[43881] + MEM[43964];
assign MEM[46874] = MEM[43882] + MEM[43972];
assign MEM[46875] = MEM[43883] + MEM[43947];
assign MEM[46876] = MEM[43885] + MEM[43958];
assign MEM[46877] = MEM[43886] + MEM[43934];
assign MEM[46878] = MEM[43887] + MEM[43930];
assign MEM[46879] = MEM[43888] + MEM[43937];
assign MEM[46880] = MEM[43889] + MEM[43965];
assign MEM[46881] = MEM[43890] + MEM[43933];
assign MEM[46882] = MEM[43891] + MEM[43936];
assign MEM[46883] = MEM[43892] + MEM[43984];
assign MEM[46884] = MEM[43896] + MEM[44008];
assign MEM[46885] = MEM[43902] + MEM[43948];
assign MEM[46886] = MEM[43903] + MEM[43932];
assign MEM[46887] = MEM[43904] + MEM[43957];
assign MEM[46888] = MEM[43905] + MEM[44011];
assign MEM[46889] = MEM[43907] + MEM[43926];
assign MEM[46890] = MEM[43908] + MEM[43968];
assign MEM[46891] = MEM[43909] + MEM[43980];
assign MEM[46892] = MEM[43910] + MEM[44015];
assign MEM[46893] = MEM[43916] + MEM[43963];
assign MEM[46894] = MEM[43918] + MEM[43949];
assign MEM[46895] = MEM[43923] + MEM[44017];
assign MEM[46896] = MEM[43924] + MEM[43971];
assign MEM[46897] = MEM[43928] + MEM[43998];
assign MEM[46898] = MEM[43931] + MEM[44012];
assign MEM[46899] = MEM[43935] + MEM[43993];
assign MEM[46900] = MEM[43938] + MEM[43990];
assign MEM[46901] = MEM[43939] + MEM[43994];
assign MEM[46902] = MEM[43940] + MEM[43985];
assign MEM[46903] = MEM[43943] + MEM[43997];
assign MEM[46904] = MEM[43944] + MEM[43983];
assign MEM[46905] = MEM[43945] + MEM[44050];
assign MEM[46906] = MEM[43946] + MEM[44004];
assign MEM[46907] = MEM[43951] + MEM[44024];
assign MEM[46908] = MEM[43952] + MEM[44005];
assign MEM[46909] = MEM[43954] + MEM[43989];
assign MEM[46910] = MEM[43955] + MEM[44029];
assign MEM[46911] = MEM[43959] + MEM[43992];
assign MEM[46912] = MEM[43960] + MEM[44000];
assign MEM[46913] = MEM[43961] + MEM[44001];
assign MEM[46914] = MEM[43962] + MEM[44006];
assign MEM[46915] = MEM[43966] + MEM[44079];
assign MEM[46916] = MEM[43967] + MEM[44014];
assign MEM[46917] = MEM[43969] + MEM[44053];
assign MEM[46918] = MEM[43973] + MEM[43991];
assign MEM[46919] = MEM[43974] + MEM[44010];
assign MEM[46920] = MEM[43975] + MEM[44021];
assign MEM[46921] = MEM[43976] + MEM[44064];
assign MEM[46922] = MEM[43977] + MEM[44054];
assign MEM[46923] = MEM[43978] + MEM[44075];
assign MEM[46924] = MEM[43979] + MEM[44052];
assign MEM[46925] = MEM[43981] + MEM[44031];
assign MEM[46926] = MEM[43982] + MEM[44055];
assign MEM[46927] = MEM[43986] + MEM[44058];
assign MEM[46928] = MEM[43988] + MEM[44087];
assign MEM[46929] = MEM[43995] + MEM[44088];
assign MEM[46930] = MEM[43996] + MEM[44030];
assign MEM[46931] = MEM[43999] + MEM[44047];
assign MEM[46932] = MEM[44002] + MEM[44091];
assign MEM[46933] = MEM[44003] + MEM[44059];
assign MEM[46934] = MEM[44007] + MEM[44038];
assign MEM[46935] = MEM[44009] + MEM[44074];
assign MEM[46936] = MEM[44013] + MEM[44063];
assign MEM[46937] = MEM[44016] + MEM[44077];
assign MEM[46938] = MEM[44018] + MEM[44107];
assign MEM[46939] = MEM[44019] + MEM[44056];
assign MEM[46940] = MEM[44020] + MEM[44073];
assign MEM[46941] = MEM[44022] + MEM[44076];
assign MEM[46942] = MEM[44023] + MEM[44112];
assign MEM[46943] = MEM[44025] + MEM[44083];
assign MEM[46944] = MEM[44026] + MEM[44118];
assign MEM[46945] = MEM[44027] + MEM[44172];
assign MEM[46946] = MEM[44028] + MEM[44126];
assign MEM[46947] = MEM[44032] + MEM[44071];
assign MEM[46948] = MEM[44033] + MEM[44143];
assign MEM[46949] = MEM[44034] + MEM[44095];
assign MEM[46950] = MEM[44035] + MEM[44096];
assign MEM[46951] = MEM[44036] + MEM[44078];
assign MEM[46952] = MEM[44037] + MEM[44108];
assign MEM[46953] = MEM[44039] + MEM[44081];
assign MEM[46954] = MEM[44040] + MEM[44110];
assign MEM[46955] = MEM[44041] + MEM[44103];
assign MEM[46956] = MEM[44042] + MEM[44105];
assign MEM[46957] = MEM[44043] + MEM[44149];
assign MEM[46958] = MEM[44044] + MEM[44089];
assign MEM[46959] = MEM[44045] + MEM[44123];
assign MEM[46960] = MEM[44046] + MEM[44099];
assign MEM[46961] = MEM[44048] + MEM[44231];
assign MEM[46962] = MEM[44049] + MEM[44145];
assign MEM[46963] = MEM[44051] + MEM[44104];
assign MEM[46964] = MEM[44057] + MEM[44125];
assign MEM[46965] = MEM[44060] + MEM[44131];
assign MEM[46966] = MEM[44061] + MEM[44148];
assign MEM[46967] = MEM[44062] + MEM[44090];
assign MEM[46968] = MEM[44065] + MEM[44214];
assign MEM[46969] = MEM[44066] + MEM[44124];
assign MEM[46970] = MEM[44067] + MEM[44102];
assign MEM[46971] = MEM[44068] + MEM[44106];
assign MEM[46972] = MEM[44069] + MEM[44162];
assign MEM[46973] = MEM[44070] + MEM[44109];
assign MEM[46974] = MEM[44072] + MEM[44139];
assign MEM[46975] = MEM[44080] + MEM[44189];
assign MEM[46976] = MEM[44082] + MEM[44156];
assign MEM[46977] = MEM[44084] + MEM[44216];
assign MEM[46978] = MEM[44085] + MEM[44163];
assign MEM[46979] = MEM[44086] + MEM[44142];
assign MEM[46980] = MEM[44092] + MEM[44136];
assign MEM[46981] = MEM[44093] + MEM[44159];
assign MEM[46982] = MEM[44094] + MEM[44169];
assign MEM[46983] = MEM[44097] + MEM[44182];
assign MEM[46984] = MEM[44098] + MEM[44161];
assign MEM[46985] = MEM[44100] + MEM[44211];
assign MEM[46986] = MEM[44101] + MEM[44166];
assign MEM[46987] = MEM[44111] + MEM[44146];
assign MEM[46988] = MEM[44113] + MEM[44160];
assign MEM[46989] = MEM[44114] + MEM[44151];
assign MEM[46990] = MEM[44115] + MEM[44128];
assign MEM[46991] = MEM[44116] + MEM[44179];
assign MEM[46992] = MEM[44117] + MEM[44173];
assign MEM[46993] = MEM[44119] + MEM[44193];
assign MEM[46994] = MEM[44120] + MEM[44209];
assign MEM[46995] = MEM[44121] + MEM[44157];
assign MEM[46996] = MEM[44122] + MEM[44165];
assign MEM[46997] = MEM[44127] + MEM[44203];
assign MEM[46998] = MEM[44129] + MEM[44212];
assign MEM[46999] = MEM[44130] + MEM[44176];
assign MEM[47000] = MEM[44132] + MEM[44178];
assign MEM[47001] = MEM[44133] + MEM[44205];
assign MEM[47002] = MEM[44134] + MEM[44191];
assign MEM[47003] = MEM[44135] + MEM[44232];
assign MEM[47004] = MEM[44137] + MEM[44184];
assign MEM[47005] = MEM[44138] + MEM[44218];
assign MEM[47006] = MEM[44140] + MEM[44217];
assign MEM[47007] = MEM[44141] + MEM[44194];
assign MEM[47008] = MEM[44144] + MEM[44196];
assign MEM[47009] = MEM[44147] + MEM[44206];
assign MEM[47010] = MEM[44150] + MEM[44195];
assign MEM[47011] = MEM[44152] + MEM[44226];
assign MEM[47012] = MEM[44153] + MEM[44188];
assign MEM[47013] = MEM[44154] + MEM[44220];
assign MEM[47014] = MEM[44155] + MEM[44202];
assign MEM[47015] = MEM[44158] + MEM[44223];
assign MEM[47016] = MEM[44164] + MEM[44222];
assign MEM[47017] = MEM[44167] + MEM[44272];
assign MEM[47018] = MEM[44168] + MEM[44239];
assign MEM[47019] = MEM[44170] + MEM[44280];
assign MEM[47020] = MEM[44171] + MEM[44198];
assign MEM[47021] = MEM[44174] + MEM[44227];
assign MEM[47022] = MEM[44175] + MEM[44215];
assign MEM[47023] = MEM[44177] + MEM[44259];
assign MEM[47024] = MEM[44180] + MEM[44299];
assign MEM[47025] = MEM[44181] + MEM[44268];
assign MEM[47026] = MEM[44183] + MEM[44251];
assign MEM[47027] = MEM[44185] + MEM[44271];
assign MEM[47028] = MEM[44186] + MEM[44240];
assign MEM[47029] = MEM[44187] + MEM[44308];
assign MEM[47030] = MEM[44190] + MEM[44267];
assign MEM[47031] = MEM[44192] + MEM[44273];
assign MEM[47032] = MEM[44197] + MEM[44322];
assign MEM[47033] = MEM[44199] + MEM[44317];
assign MEM[47034] = MEM[44200] + MEM[44287];
assign MEM[47035] = MEM[44201] + MEM[44260];
assign MEM[47036] = MEM[44204] + MEM[44295];
assign MEM[47037] = MEM[44207] + MEM[44250];
assign MEM[47038] = MEM[44208] + MEM[44291];
assign MEM[47039] = MEM[44210] + MEM[44233];
assign MEM[47040] = MEM[44213] + MEM[44241];
assign MEM[47041] = MEM[44219] + MEM[44263];
assign MEM[47042] = MEM[44221] + MEM[44245];
assign MEM[47043] = MEM[44224] + MEM[44296];
assign MEM[47044] = MEM[44225] + MEM[44278];
assign MEM[47045] = MEM[44228] + MEM[44294];
assign MEM[47046] = MEM[44229] + MEM[44325];
assign MEM[47047] = MEM[44230] + MEM[44247];
assign MEM[47048] = MEM[44234] + MEM[44289];
assign MEM[47049] = MEM[44235] + MEM[44277];
assign MEM[47050] = MEM[44236] + MEM[44284];
assign MEM[47051] = MEM[44237] + MEM[44297];
assign MEM[47052] = MEM[44238] + MEM[44281];
assign MEM[47053] = MEM[44242] + MEM[44330];
assign MEM[47054] = MEM[44243] + MEM[44275];
assign MEM[47055] = MEM[44244] + MEM[44313];
assign MEM[47056] = MEM[44246] + MEM[44293];
assign MEM[47057] = MEM[44248] + MEM[44378];
assign MEM[47058] = MEM[44249] + MEM[44333];
assign MEM[47059] = MEM[44252] + MEM[44286];
assign MEM[47060] = MEM[44253] + MEM[44318];
assign MEM[47061] = MEM[44254] + MEM[44359];
assign MEM[47062] = MEM[44255] + MEM[44298];
assign MEM[47063] = MEM[44256] + MEM[44341];
assign MEM[47064] = MEM[44257] + MEM[44315];
assign MEM[47065] = MEM[44258] + MEM[44332];
assign MEM[47066] = MEM[44261] + MEM[44303];
assign MEM[47067] = MEM[44262] + MEM[44438];
assign MEM[47068] = MEM[44264] + MEM[44405];
assign MEM[47069] = MEM[44265] + MEM[44306];
assign MEM[47070] = MEM[44266] + MEM[44336];
assign MEM[47071] = MEM[44269] + MEM[44362];
assign MEM[47072] = MEM[44270] + MEM[44312];
assign MEM[47073] = MEM[44274] + MEM[44307];
assign MEM[47074] = MEM[44276] + MEM[44329];
assign MEM[47075] = MEM[44279] + MEM[44395];
assign MEM[47076] = MEM[44282] + MEM[44413];
assign MEM[47077] = MEM[44283] + MEM[44390];
assign MEM[47078] = MEM[44285] + MEM[44335];
assign MEM[47079] = MEM[44288] + MEM[44401];
assign MEM[47080] = MEM[44290] + MEM[44348];
assign MEM[47081] = MEM[44292] + MEM[44392];
assign MEM[47082] = MEM[44300] + MEM[44327];
assign MEM[47083] = MEM[44301] + MEM[44387];
assign MEM[47084] = MEM[44302] + MEM[44337];
assign MEM[47085] = MEM[44304] + MEM[44381];
assign MEM[47086] = MEM[44305] + MEM[44463];
assign MEM[47087] = MEM[44309] + MEM[44408];
assign MEM[47088] = MEM[44310] + MEM[44376];
assign MEM[47089] = MEM[44311] + MEM[44356];
assign MEM[47090] = MEM[44314] + MEM[44345];
assign MEM[47091] = MEM[44316] + MEM[44367];
assign MEM[47092] = MEM[44319] + MEM[44361];
assign MEM[47093] = MEM[44320] + MEM[44396];
assign MEM[47094] = MEM[44321] + MEM[44377];
assign MEM[47095] = MEM[44323] + MEM[44470];
assign MEM[47096] = MEM[44324] + MEM[44353];
assign MEM[47097] = MEM[44326] + MEM[44437];
assign MEM[47098] = MEM[44328] + MEM[44372];
assign MEM[47099] = MEM[44331] + MEM[44357];
assign MEM[47100] = MEM[44334] + MEM[44399];
assign MEM[47101] = MEM[44338] + MEM[44369];
assign MEM[47102] = MEM[44339] + MEM[44363];
assign MEM[47103] = MEM[44340] + MEM[44383];
assign MEM[47104] = MEM[44342] + MEM[44404];
assign MEM[47105] = MEM[44343] + MEM[44453];
assign MEM[47106] = MEM[44344] + MEM[44393];
assign MEM[47107] = MEM[44346] + MEM[44427];
assign MEM[47108] = MEM[44347] + MEM[44474];
assign MEM[47109] = MEM[44349] + MEM[44436];
assign MEM[47110] = MEM[44350] + MEM[44384];
assign MEM[47111] = MEM[44351] + MEM[44449];
assign MEM[47112] = MEM[44352] + MEM[44366];
assign MEM[47113] = MEM[44354] + MEM[44410];
assign MEM[47114] = MEM[44355] + MEM[44388];
assign MEM[47115] = MEM[44358] + MEM[44426];
assign MEM[47116] = MEM[44360] + MEM[44412];
assign MEM[47117] = MEM[44364] + MEM[44403];
assign MEM[47118] = MEM[44365] + MEM[44503];
assign MEM[47119] = MEM[44368] + MEM[44418];
assign MEM[47120] = MEM[44370] + MEM[44421];
assign MEM[47121] = MEM[44371] + MEM[44406];
assign MEM[47122] = MEM[44373] + MEM[44429];
assign MEM[47123] = MEM[44374] + MEM[44409];
assign MEM[47124] = MEM[44375] + MEM[44423];
assign MEM[47125] = MEM[44379] + MEM[44516];
assign MEM[47126] = MEM[44380] + MEM[44398];
assign MEM[47127] = MEM[44382] + MEM[44428];
assign MEM[47128] = MEM[44385] + MEM[44435];
assign MEM[47129] = MEM[44386] + MEM[44496];
assign MEM[47130] = MEM[44389] + MEM[44459];
assign MEM[47131] = MEM[44391] + MEM[44424];
assign MEM[47132] = MEM[44394] + MEM[44486];
assign MEM[47133] = MEM[44397] + MEM[44460];
assign MEM[47134] = MEM[44400] + MEM[44443];
assign MEM[47135] = MEM[44402] + MEM[44444];
assign MEM[47136] = MEM[44407] + MEM[44483];
assign MEM[47137] = MEM[44411] + MEM[44446];
assign MEM[47138] = MEM[44414] + MEM[44484];
assign MEM[47139] = MEM[44415] + MEM[44473];
assign MEM[47140] = MEM[44416] + MEM[44471];
assign MEM[47141] = MEM[44417] + MEM[44456];
assign MEM[47142] = MEM[44419] + MEM[44442];
assign MEM[47143] = MEM[44420] + MEM[44454];
assign MEM[47144] = MEM[44422] + MEM[44455];
assign MEM[47145] = MEM[44425] + MEM[44491];
assign MEM[47146] = MEM[44430] + MEM[44494];
assign MEM[47147] = MEM[44431] + MEM[44552];
assign MEM[47148] = MEM[44432] + MEM[44506];
assign MEM[47149] = MEM[44433] + MEM[44517];
assign MEM[47150] = MEM[44434] + MEM[44477];
assign MEM[47151] = MEM[44439] + MEM[44553];
assign MEM[47152] = MEM[44440] + MEM[44505];
assign MEM[47153] = MEM[44441] + MEM[44580];
assign MEM[47154] = MEM[44445] + MEM[44504];
assign MEM[47155] = MEM[44447] + MEM[44476];
assign MEM[47156] = MEM[44448] + MEM[44489];
assign MEM[47157] = MEM[44450] + MEM[44520];
assign MEM[47158] = MEM[44451] + MEM[44540];
assign MEM[47159] = MEM[44452] + MEM[44582];
assign MEM[47160] = MEM[44457] + MEM[44524];
assign MEM[47161] = MEM[44458] + MEM[44523];
assign MEM[47162] = MEM[44461] + MEM[44555];
assign MEM[47163] = MEM[44462] + MEM[44507];
assign MEM[47164] = MEM[44464] + MEM[44533];
assign MEM[47165] = MEM[44465] + MEM[44525];
assign MEM[47166] = MEM[44466] + MEM[44548];
assign MEM[47167] = MEM[44467] + MEM[44513];
assign MEM[47168] = MEM[44468] + MEM[44508];
assign MEM[47169] = MEM[44469] + MEM[44536];
assign MEM[47170] = MEM[44472] + MEM[44539];
assign MEM[47171] = MEM[44475] + MEM[44511];
assign MEM[47172] = MEM[44478] + MEM[44502];
assign MEM[47173] = MEM[44479] + MEM[44574];
assign MEM[47174] = MEM[44480] + MEM[44530];
assign MEM[47175] = MEM[44481] + MEM[44542];
assign MEM[47176] = MEM[44482] + MEM[44638];
assign MEM[47177] = MEM[44485] + MEM[44537];
assign MEM[47178] = MEM[44487] + MEM[44550];
assign MEM[47179] = MEM[44488] + MEM[44576];
assign MEM[47180] = MEM[44490] + MEM[44560];
assign MEM[47181] = MEM[44492] + MEM[44586];
assign MEM[47182] = MEM[44493] + MEM[44534];
assign MEM[47183] = MEM[44495] + MEM[44529];
assign MEM[47184] = MEM[44497] + MEM[44572];
assign MEM[47185] = MEM[44498] + MEM[44570];
assign MEM[47186] = MEM[44499] + MEM[44531];
assign MEM[47187] = MEM[44500] + MEM[44604];
assign MEM[47188] = MEM[44501] + MEM[44623];
assign MEM[47189] = MEM[44509] + MEM[44554];
assign MEM[47190] = MEM[44510] + MEM[44577];
assign MEM[47191] = MEM[44512] + MEM[44535];
assign MEM[47192] = MEM[44514] + MEM[44607];
assign MEM[47193] = MEM[44515] + MEM[44588];
assign MEM[47194] = MEM[44518] + MEM[44625];
assign MEM[47195] = MEM[44519] + MEM[44589];
assign MEM[47196] = MEM[44521] + MEM[44611];
assign MEM[47197] = MEM[44522] + MEM[44606];
assign MEM[47198] = MEM[44526] + MEM[44600];
assign MEM[47199] = MEM[44527] + MEM[44559];
assign MEM[47200] = MEM[44528] + MEM[44624];
assign MEM[47201] = MEM[44532] + MEM[44557];
assign MEM[47202] = MEM[44538] + MEM[44601];
assign MEM[47203] = MEM[44541] + MEM[44617];
assign MEM[47204] = MEM[44543] + MEM[44614];
assign MEM[47205] = MEM[44544] + MEM[44621];
assign MEM[47206] = MEM[44545] + MEM[44571];
assign MEM[47207] = MEM[44546] + MEM[44696];
assign MEM[47208] = MEM[44547] + MEM[44605];
assign MEM[47209] = MEM[44549] + MEM[44642];
assign MEM[47210] = MEM[44551] + MEM[44630];
assign MEM[47211] = MEM[44556] + MEM[44569];
assign MEM[47212] = MEM[44558] + MEM[44662];
assign MEM[47213] = MEM[44561] + MEM[44629];
assign MEM[47214] = MEM[44562] + MEM[44669];
assign MEM[47215] = MEM[44563] + MEM[44655];
assign MEM[47216] = MEM[44564] + MEM[44595];
assign MEM[47217] = MEM[44565] + MEM[44616];
assign MEM[47218] = MEM[44566] + MEM[44690];
assign MEM[47219] = MEM[44567] + MEM[44631];
assign MEM[47220] = MEM[44568] + MEM[44639];
assign MEM[47221] = MEM[44573] + MEM[44599];
assign MEM[47222] = MEM[44575] + MEM[44646];
assign MEM[47223] = MEM[44578] + MEM[44626];
assign MEM[47224] = MEM[44579] + MEM[44636];
assign MEM[47225] = MEM[44581] + MEM[44660];
assign MEM[47226] = MEM[44583] + MEM[44613];
assign MEM[47227] = MEM[44584] + MEM[44680];
assign MEM[47228] = MEM[44585] + MEM[44674];
assign MEM[47229] = MEM[44587] + MEM[44633];
assign MEM[47230] = MEM[44590] + MEM[44648];
assign MEM[47231] = MEM[44591] + MEM[44615];
assign MEM[47232] = MEM[44592] + MEM[44667];
assign MEM[47233] = MEM[44593] + MEM[44628];
assign MEM[47234] = MEM[44594] + MEM[44657];
assign MEM[47235] = MEM[44596] + MEM[44643];
assign MEM[47236] = MEM[44597] + MEM[44730];
assign MEM[47237] = MEM[44598] + MEM[44640];
assign MEM[47238] = MEM[44602] + MEM[44649];
assign MEM[47239] = MEM[44603] + MEM[44670];
assign MEM[47240] = MEM[44608] + MEM[44738];
assign MEM[47241] = MEM[44609] + MEM[44722];
assign MEM[47242] = MEM[44610] + MEM[44644];
assign MEM[47243] = MEM[44612] + MEM[44656];
assign MEM[47244] = MEM[44618] + MEM[44678];
assign MEM[47245] = MEM[44619] + MEM[44651];
assign MEM[47246] = MEM[44620] + MEM[44677];
assign MEM[47247] = MEM[44622] + MEM[44652];
assign MEM[47248] = MEM[44627] + MEM[44675];
assign MEM[47249] = MEM[44632] + MEM[44712];
assign MEM[47250] = MEM[44634] + MEM[44704];
assign MEM[47251] = MEM[44635] + MEM[44701];
assign MEM[47252] = MEM[44637] + MEM[44747];
assign MEM[47253] = MEM[44641] + MEM[44686];
assign MEM[47254] = MEM[44645] + MEM[44709];
assign MEM[47255] = MEM[44647] + MEM[44723];
assign MEM[47256] = MEM[44650] + MEM[44697];
assign MEM[47257] = MEM[44653] + MEM[44689];
assign MEM[47258] = MEM[44654] + MEM[44707];
assign MEM[47259] = MEM[44658] + MEM[44753];
assign MEM[47260] = MEM[44659] + MEM[44756];
assign MEM[47261] = MEM[44661] + MEM[44732];
assign MEM[47262] = MEM[44663] + MEM[44692];
assign MEM[47263] = MEM[44664] + MEM[44706];
assign MEM[47264] = MEM[44665] + MEM[44758];
assign MEM[47265] = MEM[44666] + MEM[44744];
assign MEM[47266] = MEM[44668] + MEM[44694];
assign MEM[47267] = MEM[44671] + MEM[44780];
assign MEM[47268] = MEM[44672] + MEM[44728];
assign MEM[47269] = MEM[44673] + MEM[44798];
assign MEM[47270] = MEM[44676] + MEM[44731];
assign MEM[47271] = MEM[44679] + MEM[44789];
assign MEM[47272] = MEM[44681] + MEM[44715];
assign MEM[47273] = MEM[44682] + MEM[44762];
assign MEM[47274] = MEM[44683] + MEM[44725];
assign MEM[47275] = MEM[44684] + MEM[44736];
assign MEM[47276] = MEM[44685] + MEM[44766];
assign MEM[47277] = MEM[44687] + MEM[44792];
assign MEM[47278] = MEM[44688] + MEM[44757];
assign MEM[47279] = MEM[44691] + MEM[44783];
assign MEM[47280] = MEM[44693] + MEM[44743];
assign MEM[47281] = MEM[44695] + MEM[44750];
assign MEM[47282] = MEM[44698] + MEM[44781];
assign MEM[47283] = MEM[44699] + MEM[44735];
assign MEM[47284] = MEM[44700] + MEM[44835];
assign MEM[47285] = MEM[44702] + MEM[44803];
assign MEM[47286] = MEM[44703] + MEM[44729];
assign MEM[47287] = MEM[44705] + MEM[44791];
assign MEM[47288] = MEM[44708] + MEM[44734];
assign MEM[47289] = MEM[44710] + MEM[44839];
assign MEM[47290] = MEM[44711] + MEM[44749];
assign MEM[47291] = MEM[44713] + MEM[44802];
assign MEM[47292] = MEM[44714] + MEM[44778];
assign MEM[47293] = MEM[44716] + MEM[44824];
assign MEM[47294] = MEM[44717] + MEM[44740];
assign MEM[47295] = MEM[44718] + MEM[44777];
assign MEM[47296] = MEM[44719] + MEM[44813];
assign MEM[47297] = MEM[44720] + MEM[44771];
assign MEM[47298] = MEM[44721] + MEM[44814];
assign MEM[47299] = MEM[44724] + MEM[44755];
assign MEM[47300] = MEM[44726] + MEM[44745];
assign MEM[47301] = MEM[44727] + MEM[44795];
assign MEM[47302] = MEM[44733] + MEM[44770];
assign MEM[47303] = MEM[44737] + MEM[44806];
assign MEM[47304] = MEM[44739] + MEM[44764];
assign MEM[47305] = MEM[44741] + MEM[44793];
assign MEM[47306] = MEM[44742] + MEM[44784];
assign MEM[47307] = MEM[44746] + MEM[44774];
assign MEM[47308] = MEM[44748] + MEM[44843];
assign MEM[47309] = MEM[44751] + MEM[44818];
assign MEM[47310] = MEM[44752] + MEM[44828];
assign MEM[47311] = MEM[44754] + MEM[44858];
assign MEM[47312] = MEM[44759] + MEM[44845];
assign MEM[47313] = MEM[44760] + MEM[44815];
assign MEM[47314] = MEM[44761] + MEM[44825];
assign MEM[47315] = MEM[44763] + MEM[44801];
assign MEM[47316] = MEM[44765] + MEM[44810];
assign MEM[47317] = MEM[44767] + MEM[44836];
assign MEM[47318] = MEM[44768] + MEM[44811];
assign MEM[47319] = MEM[44769] + MEM[44809];
assign MEM[47320] = MEM[44772] + MEM[44855];
assign MEM[47321] = MEM[44773] + MEM[44788];
assign MEM[47322] = MEM[44775] + MEM[44863];
assign MEM[47323] = MEM[44776] + MEM[44850];
assign MEM[47324] = MEM[44779] + MEM[44867];
assign MEM[47325] = MEM[44782] + MEM[44906];
assign MEM[47326] = MEM[44785] + MEM[44967];
assign MEM[47327] = MEM[44786] + MEM[44807];
assign MEM[47328] = MEM[44787] + MEM[44859];
assign MEM[47329] = MEM[44790] + MEM[44817];
assign MEM[47330] = MEM[44794] + MEM[44805];
assign MEM[47331] = MEM[44796] + MEM[44865];
assign MEM[47332] = MEM[44797] + MEM[44864];
assign MEM[47333] = MEM[44799] + MEM[44854];
assign MEM[47334] = MEM[44800] + MEM[44861];
assign MEM[47335] = MEM[44804] + MEM[44866];
assign MEM[47336] = MEM[44808] + MEM[44885];
assign MEM[47337] = MEM[44812] + MEM[44900];
assign MEM[47338] = MEM[44816] + MEM[44884];
assign MEM[47339] = MEM[44819] + MEM[44860];
assign MEM[47340] = MEM[44820] + MEM[44938];
assign MEM[47341] = MEM[44821] + MEM[44876];
assign MEM[47342] = MEM[44822] + MEM[44862];
assign MEM[47343] = MEM[44823] + MEM[44880];
assign MEM[47344] = MEM[44826] + MEM[44878];
assign MEM[47345] = MEM[44827] + MEM[44870];
assign MEM[47346] = MEM[44829] + MEM[44851];
assign MEM[47347] = MEM[44830] + MEM[44890];
assign MEM[47348] = MEM[44831] + MEM[44888];
assign MEM[47349] = MEM[44832] + MEM[44872];
assign MEM[47350] = MEM[44833] + MEM[44904];
assign MEM[47351] = MEM[44834] + MEM[44853];
assign MEM[47352] = MEM[44837] + MEM[44868];
assign MEM[47353] = MEM[44838] + MEM[44891];
assign MEM[47354] = MEM[44840] + MEM[44970];
assign MEM[47355] = MEM[44841] + MEM[44952];
assign MEM[47356] = MEM[44842] + MEM[44902];
assign MEM[47357] = MEM[44844] + MEM[44897];
assign MEM[47358] = MEM[44846] + MEM[44887];
assign MEM[47359] = MEM[44847] + MEM[45022];
assign MEM[47360] = MEM[44848] + MEM[44939];
assign MEM[47361] = MEM[44849] + MEM[44881];
assign MEM[47362] = MEM[44852] + MEM[45016];
assign MEM[47363] = MEM[44856] + MEM[44931];
assign MEM[47364] = MEM[44857] + MEM[44886];
assign MEM[47365] = MEM[44869] + MEM[44932];
assign MEM[47366] = MEM[44871] + MEM[44909];
assign MEM[47367] = MEM[44873] + MEM[44943];
assign MEM[47368] = MEM[44874] + MEM[44935];
assign MEM[47369] = MEM[44875] + MEM[44942];
assign MEM[47370] = MEM[44877] + MEM[44977];
assign MEM[47371] = MEM[44879] + MEM[44922];
assign MEM[47372] = MEM[44882] + MEM[44915];
assign MEM[47373] = MEM[44883] + MEM[44960];
assign MEM[47374] = MEM[44889] + MEM[44995];
assign MEM[47375] = MEM[44892] + MEM[44930];
assign MEM[47376] = MEM[44893] + MEM[44936];
assign MEM[47377] = MEM[44894] + MEM[44969];
assign MEM[47378] = MEM[44895] + MEM[45011];
assign MEM[47379] = MEM[44896] + MEM[44997];
assign MEM[47380] = MEM[44898] + MEM[44933];
assign MEM[47381] = MEM[44899] + MEM[44907];
assign MEM[47382] = MEM[44901] + MEM[44966];
assign MEM[47383] = MEM[44903] + MEM[44946];
assign MEM[47384] = MEM[44905] + MEM[44965];
assign MEM[47385] = MEM[44908] + MEM[44973];
assign MEM[47386] = MEM[44910] + MEM[45001];
assign MEM[47387] = MEM[44911] + MEM[44964];
assign MEM[47388] = MEM[44912] + MEM[45014];
assign MEM[47389] = MEM[44913] + MEM[44949];
assign MEM[47390] = MEM[44914] + MEM[45002];
assign MEM[47391] = MEM[44916] + MEM[45010];
assign MEM[47392] = MEM[44917] + MEM[45009];
assign MEM[47393] = MEM[44918] + MEM[44951];
assign MEM[47394] = MEM[44919] + MEM[44954];
assign MEM[47395] = MEM[44920] + MEM[44959];
assign MEM[47396] = MEM[44921] + MEM[44955];
assign MEM[47397] = MEM[44923] + MEM[45000];
assign MEM[47398] = MEM[44924] + MEM[44986];
assign MEM[47399] = MEM[44925] + MEM[44974];
assign MEM[47400] = MEM[44926] + MEM[45005];
assign MEM[47401] = MEM[44927] + MEM[44993];
assign MEM[47402] = MEM[44928] + MEM[44990];
assign MEM[47403] = MEM[44929] + MEM[44957];
assign MEM[47404] = MEM[44934] + MEM[45037];
assign MEM[47405] = MEM[44937] + MEM[45030];
assign MEM[47406] = MEM[44940] + MEM[44981];
assign MEM[47407] = MEM[44941] + MEM[44984];
assign MEM[47408] = MEM[44944] + MEM[44976];
assign MEM[47409] = MEM[44945] + MEM[44962];
assign MEM[47410] = MEM[44947] + MEM[45055];
assign MEM[47411] = MEM[44948] + MEM[45046];
assign MEM[47412] = MEM[44950] + MEM[45031];
assign MEM[47413] = MEM[44953] + MEM[44987];
assign MEM[47414] = MEM[44956] + MEM[45039];
assign MEM[47415] = MEM[44958] + MEM[45034];
assign MEM[47416] = MEM[44961] + MEM[44983];
assign MEM[47417] = MEM[44963] + MEM[45013];
assign MEM[47418] = MEM[44968] + MEM[44992];
assign MEM[47419] = MEM[44971] + MEM[45015];
assign MEM[47420] = MEM[44972] + MEM[45019];
assign MEM[47421] = MEM[44975] + MEM[45021];
assign MEM[47422] = MEM[44978] + MEM[45012];
assign MEM[47423] = MEM[44979] + MEM[45057];
assign MEM[47424] = MEM[44980] + MEM[45024];
assign MEM[47425] = MEM[44982] + MEM[45091];
assign MEM[47426] = MEM[44985] + MEM[45062];
assign MEM[47427] = MEM[44988] + MEM[45064];
assign MEM[47428] = MEM[44989] + MEM[45061];
assign MEM[47429] = MEM[44991] + MEM[45144];
assign MEM[47430] = MEM[44994] + MEM[45056];
assign MEM[47431] = MEM[44996] + MEM[45115];
assign MEM[47432] = MEM[44998] + MEM[45047];
assign MEM[47433] = MEM[44999] + MEM[45027];
assign MEM[47434] = MEM[45003] + MEM[45095];
assign MEM[47435] = MEM[45004] + MEM[45086];
assign MEM[47436] = MEM[45006] + MEM[45040];
assign MEM[47437] = MEM[45007] + MEM[45075];
assign MEM[47438] = MEM[45008] + MEM[45051];
assign MEM[47439] = MEM[45017] + MEM[45104];
assign MEM[47440] = MEM[45018] + MEM[45139];
assign MEM[47441] = MEM[45020] + MEM[45054];
assign MEM[47442] = MEM[45023] + MEM[45090];
assign MEM[47443] = MEM[45025] + MEM[45082];
assign MEM[47444] = MEM[45026] + MEM[45074];
assign MEM[47445] = MEM[45028] + MEM[45078];
assign MEM[47446] = MEM[45029] + MEM[45080];
assign MEM[47447] = MEM[45032] + MEM[45058];
assign MEM[47448] = MEM[45033] + MEM[45140];
assign MEM[47449] = MEM[45035] + MEM[45094];
assign MEM[47450] = MEM[45036] + MEM[45112];
assign MEM[47451] = MEM[45038] + MEM[45084];
assign MEM[47452] = MEM[45041] + MEM[45118];
assign MEM[47453] = MEM[45042] + MEM[45123];
assign MEM[47454] = MEM[45043] + MEM[45079];
assign MEM[47455] = MEM[45044] + MEM[45108];
assign MEM[47456] = MEM[45045] + MEM[45076];
assign MEM[47457] = MEM[45048] + MEM[45093];
assign MEM[47458] = MEM[45049] + MEM[45083];
assign MEM[47459] = MEM[45050] + MEM[45138];
assign MEM[47460] = MEM[45052] + MEM[45125];
assign MEM[47461] = MEM[45053] + MEM[45128];
assign MEM[47462] = MEM[45059] + MEM[45087];
assign MEM[47463] = MEM[45060] + MEM[45096];
assign MEM[47464] = MEM[45063] + MEM[45122];
assign MEM[47465] = MEM[45065] + MEM[45178];
assign MEM[47466] = MEM[45066] + MEM[45111];
assign MEM[47467] = MEM[45067] + MEM[45147];
assign MEM[47468] = MEM[45068] + MEM[45135];
assign MEM[47469] = MEM[45069] + MEM[45145];
assign MEM[47470] = MEM[45070] + MEM[45097];
assign MEM[47471] = MEM[45071] + MEM[45168];
assign MEM[47472] = MEM[45072] + MEM[45166];
assign MEM[47473] = MEM[45073] + MEM[45132];
assign MEM[47474] = MEM[45077] + MEM[45154];
assign MEM[47475] = MEM[45081] + MEM[45167];
assign MEM[47476] = MEM[45085] + MEM[45155];
assign MEM[47477] = MEM[45088] + MEM[45186];
assign MEM[47478] = MEM[45089] + MEM[45171];
assign MEM[47479] = MEM[45092] + MEM[45106];
assign MEM[47480] = MEM[45098] + MEM[45148];
assign MEM[47481] = MEM[45099] + MEM[45193];
assign MEM[47482] = MEM[45100] + MEM[45151];
assign MEM[47483] = MEM[45101] + MEM[45153];
assign MEM[47484] = MEM[45102] + MEM[45157];
assign MEM[47485] = MEM[45103] + MEM[45172];
assign MEM[47486] = MEM[45105] + MEM[45146];
assign MEM[47487] = MEM[45107] + MEM[45127];
assign MEM[47488] = MEM[45109] + MEM[45116];
assign MEM[47489] = MEM[45110] + MEM[45182];
assign MEM[47490] = MEM[45113] + MEM[45199];
assign MEM[47491] = MEM[45114] + MEM[45185];
assign MEM[47492] = MEM[45117] + MEM[45165];
assign MEM[47493] = MEM[45119] + MEM[45179];
assign MEM[47494] = MEM[45120] + MEM[45180];
assign MEM[47495] = MEM[45121] + MEM[45203];
assign MEM[47496] = MEM[45124] + MEM[45189];
assign MEM[47497] = MEM[45126] + MEM[45175];
assign MEM[47498] = MEM[45129] + MEM[45257];
assign MEM[47499] = MEM[45130] + MEM[45174];
assign MEM[47500] = MEM[45131] + MEM[45176];
assign MEM[47501] = MEM[45133] + MEM[45233];
assign MEM[47502] = MEM[45134] + MEM[45198];
assign MEM[47503] = MEM[45136] + MEM[45194];
assign MEM[47504] = MEM[45137] + MEM[45239];
assign MEM[47505] = MEM[45141] + MEM[45160];
assign MEM[47506] = MEM[45142] + MEM[45229];
assign MEM[47507] = MEM[45143] + MEM[45208];
assign MEM[47508] = MEM[45149] + MEM[45275];
assign MEM[47509] = MEM[45150] + MEM[45183];
assign MEM[47510] = MEM[45152] + MEM[45235];
assign MEM[47511] = MEM[45156] + MEM[45223];
assign MEM[47512] = MEM[45158] + MEM[45303];
assign MEM[47513] = MEM[45159] + MEM[45216];
assign MEM[47514] = MEM[45161] + MEM[45230];
assign MEM[47515] = MEM[45162] + MEM[45249];
assign MEM[47516] = MEM[45163] + MEM[45192];
assign MEM[47517] = MEM[45164] + MEM[45205];
assign MEM[47518] = MEM[45169] + MEM[45261];
assign MEM[47519] = MEM[45170] + MEM[45244];
assign MEM[47520] = MEM[45173] + MEM[45301];
assign MEM[47521] = MEM[45177] + MEM[45236];
assign MEM[47522] = MEM[45181] + MEM[45227];
assign MEM[47523] = MEM[45184] + MEM[45209];
assign MEM[47524] = MEM[45187] + MEM[45242];
assign MEM[47525] = MEM[45188] + MEM[45302];
assign MEM[47526] = MEM[45190] + MEM[45272];
assign MEM[47527] = MEM[45191] + MEM[45283];
assign MEM[47528] = MEM[45195] + MEM[45270];
assign MEM[47529] = MEM[45196] + MEM[45251];
assign MEM[47530] = MEM[45197] + MEM[45290];
assign MEM[47531] = MEM[45200] + MEM[45245];
assign MEM[47532] = MEM[45201] + MEM[45356];
assign MEM[47533] = MEM[45202] + MEM[45259];
assign MEM[47534] = MEM[45204] + MEM[45248];
assign MEM[47535] = MEM[45206] + MEM[45264];
assign MEM[47536] = MEM[45207] + MEM[45255];
assign MEM[47537] = MEM[45210] + MEM[45241];
assign MEM[47538] = MEM[45211] + MEM[45346];
assign MEM[47539] = MEM[45212] + MEM[45265];
assign MEM[47540] = MEM[45213] + MEM[45231];
assign MEM[47541] = MEM[45214] + MEM[45350];
assign MEM[47542] = MEM[45215] + MEM[45289];
assign MEM[47543] = MEM[45217] + MEM[45305];
assign MEM[47544] = MEM[45218] + MEM[45267];
assign MEM[47545] = MEM[45219] + MEM[45291];
assign MEM[47546] = MEM[45220] + MEM[45258];
assign MEM[47547] = MEM[45221] + MEM[45297];
assign MEM[47548] = MEM[45222] + MEM[45274];
assign MEM[47549] = MEM[45224] + MEM[45252];
assign MEM[47550] = MEM[45225] + MEM[45253];
assign MEM[47551] = MEM[45226] + MEM[45263];
assign MEM[47552] = MEM[45228] + MEM[45260];
assign MEM[47553] = MEM[45232] + MEM[45324];
assign MEM[47554] = MEM[45234] + MEM[45299];
assign MEM[47555] = MEM[45237] + MEM[45317];
assign MEM[47556] = MEM[45238] + MEM[45298];
assign MEM[47557] = MEM[45240] + MEM[45287];
assign MEM[47558] = MEM[45243] + MEM[45280];
assign MEM[47559] = MEM[45246] + MEM[45304];
assign MEM[47560] = MEM[45247] + MEM[45348];
assign MEM[47561] = MEM[45250] + MEM[45329];
assign MEM[47562] = MEM[45254] + MEM[45337];
assign MEM[47563] = MEM[45256] + MEM[45322];
assign MEM[47564] = MEM[45262] + MEM[45296];
assign MEM[47565] = MEM[45266] + MEM[45334];
assign MEM[47566] = MEM[45268] + MEM[45327];
assign MEM[47567] = MEM[45269] + MEM[45320];
assign MEM[47568] = MEM[45271] + MEM[45310];
assign MEM[47569] = MEM[45273] + MEM[45377];
assign MEM[47570] = MEM[45276] + MEM[45315];
assign MEM[47571] = MEM[45277] + MEM[45319];
assign MEM[47572] = MEM[45278] + MEM[45323];
assign MEM[47573] = MEM[45279] + MEM[45331];
assign MEM[47574] = MEM[45281] + MEM[45351];
assign MEM[47575] = MEM[45282] + MEM[45366];
assign MEM[47576] = MEM[45284] + MEM[45398];
assign MEM[47577] = MEM[45285] + MEM[45345];
assign MEM[47578] = MEM[45286] + MEM[45400];
assign MEM[47579] = MEM[45288] + MEM[45382];
assign MEM[47580] = MEM[45292] + MEM[45333];
assign MEM[47581] = MEM[45293] + MEM[45362];
assign MEM[47582] = MEM[45294] + MEM[45363];
assign MEM[47583] = MEM[45295] + MEM[45355];
assign MEM[47584] = MEM[45300] + MEM[45376];
assign MEM[47585] = MEM[45306] + MEM[45318];
assign MEM[47586] = MEM[45307] + MEM[45419];
assign MEM[47587] = MEM[45308] + MEM[45380];
assign MEM[47588] = MEM[45309] + MEM[45421];
assign MEM[47589] = MEM[45311] + MEM[45359];
assign MEM[47590] = MEM[45312] + MEM[45445];
assign MEM[47591] = MEM[45313] + MEM[45383];
assign MEM[47592] = MEM[45314] + MEM[45373];
assign MEM[47593] = MEM[45316] + MEM[45365];
assign MEM[47594] = MEM[45321] + MEM[45425];
assign MEM[47595] = MEM[45325] + MEM[45374];
assign MEM[47596] = MEM[45326] + MEM[45372];
assign MEM[47597] = MEM[45328] + MEM[45364];
assign MEM[47598] = MEM[45330] + MEM[45395];
assign MEM[47599] = MEM[45332] + MEM[45422];
assign MEM[47600] = MEM[45335] + MEM[45384];
assign MEM[47601] = MEM[45336] + MEM[45441];
assign MEM[47602] = MEM[45338] + MEM[45357];
assign MEM[47603] = MEM[45339] + MEM[45435];
assign MEM[47604] = MEM[45340] + MEM[45367];
assign MEM[47605] = MEM[45341] + MEM[45371];
assign MEM[47606] = MEM[45342] + MEM[45412];
assign MEM[47607] = MEM[45343] + MEM[45392];
assign MEM[47608] = MEM[45344] + MEM[45389];
assign MEM[47609] = MEM[45347] + MEM[45434];
assign MEM[47610] = MEM[45349] + MEM[45410];
assign MEM[47611] = MEM[45352] + MEM[45397];
assign MEM[47612] = MEM[45353] + MEM[45420];
assign MEM[47613] = MEM[45354] + MEM[45418];
assign MEM[47614] = MEM[45358] + MEM[45406];
assign MEM[47615] = MEM[45360] + MEM[45462];
assign MEM[47616] = MEM[45361] + MEM[45409];
assign MEM[47617] = MEM[45368] + MEM[45387];
assign MEM[47618] = MEM[45369] + MEM[45428];
assign MEM[47619] = MEM[45370] + MEM[45437];
assign MEM[47620] = MEM[45375] + MEM[45467];
assign MEM[47621] = MEM[45378] + MEM[45443];
assign MEM[47622] = MEM[45379] + MEM[45414];
assign MEM[47623] = MEM[45381] + MEM[45500];
assign MEM[47624] = MEM[45385] + MEM[45469];
assign MEM[47625] = MEM[45386] + MEM[45436];
assign MEM[47626] = MEM[45388] + MEM[45449];
assign MEM[47627] = MEM[45390] + MEM[45476];
assign MEM[47628] = MEM[45391] + MEM[45454];
assign MEM[47629] = MEM[45393] + MEM[45417];
assign MEM[47630] = MEM[45394] + MEM[45470];
assign MEM[47631] = MEM[45396] + MEM[45544];
assign MEM[47632] = MEM[45399] + MEM[45447];
assign MEM[47633] = MEM[45401] + MEM[45486];
assign MEM[47634] = MEM[45402] + MEM[45455];
assign MEM[47635] = MEM[45403] + MEM[45487];
assign MEM[47636] = MEM[45404] + MEM[45466];
assign MEM[47637] = MEM[45405] + MEM[45485];
assign MEM[47638] = MEM[45407] + MEM[45498];
assign MEM[47639] = MEM[45408] + MEM[45442];
assign MEM[47640] = MEM[45411] + MEM[45453];
assign MEM[47641] = MEM[45413] + MEM[45519];
assign MEM[47642] = MEM[45415] + MEM[45460];
assign MEM[47643] = MEM[45416] + MEM[45514];
assign MEM[47644] = MEM[45423] + MEM[45505];
assign MEM[47645] = MEM[45424] + MEM[45522];
assign MEM[47646] = MEM[45426] + MEM[45491];
assign MEM[47647] = MEM[45427] + MEM[45493];
assign MEM[47648] = MEM[45429] + MEM[45457];
assign MEM[47649] = MEM[45430] + MEM[45502];
assign MEM[47650] = MEM[45431] + MEM[45490];
assign MEM[47651] = MEM[45432] + MEM[45450];
assign MEM[47652] = MEM[45433] + MEM[45465];
assign MEM[47653] = MEM[45438] + MEM[45558];
assign MEM[47654] = MEM[45439] + MEM[45479];
assign MEM[47655] = MEM[45440] + MEM[45515];
assign MEM[47656] = MEM[45444] + MEM[45569];
assign MEM[47657] = MEM[45446] + MEM[45507];
assign MEM[47658] = MEM[45448] + MEM[45496];
assign MEM[47659] = MEM[45451] + MEM[45533];
assign MEM[47660] = MEM[45452] + MEM[45478];
assign MEM[47661] = MEM[45456] + MEM[45535];
assign MEM[47662] = MEM[45458] + MEM[45520];
assign MEM[47663] = MEM[45459] + MEM[45542];
assign MEM[47664] = MEM[45461] + MEM[45506];
assign MEM[47665] = MEM[45463] + MEM[45545];
assign MEM[47666] = MEM[45464] + MEM[45543];
assign MEM[47667] = MEM[45468] + MEM[45538];
assign MEM[47668] = MEM[45471] + MEM[45510];
assign MEM[47669] = MEM[45472] + MEM[45570];
assign MEM[47670] = MEM[45473] + MEM[45594];
assign MEM[47671] = MEM[45474] + MEM[45574];
assign MEM[47672] = MEM[45475] + MEM[45534];
assign MEM[47673] = MEM[45477] + MEM[45501];
assign MEM[47674] = MEM[45480] + MEM[45529];
assign MEM[47675] = MEM[45481] + MEM[45551];
assign MEM[47676] = MEM[45482] + MEM[45523];
assign MEM[47677] = MEM[45483] + MEM[45521];
assign MEM[47678] = MEM[45484] + MEM[45539];
assign MEM[47679] = MEM[45488] + MEM[45517];
assign MEM[47680] = MEM[45489] + MEM[45548];
assign MEM[47681] = MEM[45492] + MEM[45576];
assign MEM[47682] = MEM[45494] + MEM[45552];
assign MEM[47683] = MEM[45495] + MEM[45512];
assign MEM[47684] = MEM[45497] + MEM[45584];
assign MEM[47685] = MEM[45499] + MEM[45550];
assign MEM[47686] = MEM[45503] + MEM[45566];
assign MEM[47687] = MEM[45504] + MEM[45567];
assign MEM[47688] = MEM[45508] + MEM[45620];
assign MEM[47689] = MEM[45509] + MEM[45673];
assign MEM[47690] = MEM[45511] + MEM[45568];
assign MEM[47691] = MEM[45513] + MEM[45555];
assign MEM[47692] = MEM[45516] + MEM[45615];
assign MEM[47693] = MEM[45518] + MEM[45575];
assign MEM[47694] = MEM[45524] + MEM[45633];
assign MEM[47695] = MEM[45525] + MEM[45589];
assign MEM[47696] = MEM[45526] + MEM[45588];
assign MEM[47697] = MEM[45527] + MEM[45597];
assign MEM[47698] = MEM[45528] + MEM[45572];
assign MEM[47699] = MEM[45530] + MEM[45553];
assign MEM[47700] = MEM[45531] + MEM[45605];
assign MEM[47701] = MEM[45532] + MEM[45696];
assign MEM[47702] = MEM[45536] + MEM[45647];
assign MEM[47703] = MEM[45537] + MEM[45627];
assign MEM[47704] = MEM[45540] + MEM[45608];
assign MEM[47705] = MEM[45541] + MEM[45603];
assign MEM[47706] = MEM[45546] + MEM[45665];
assign MEM[47707] = MEM[45547] + MEM[45604];
assign MEM[47708] = MEM[45549] + MEM[45580];
assign MEM[47709] = MEM[45554] + MEM[45577];
assign MEM[47710] = MEM[45556] + MEM[45610];
assign MEM[47711] = MEM[45557] + MEM[45614];
assign MEM[47712] = MEM[45559] + MEM[45663];
assign MEM[47713] = MEM[45560] + MEM[45613];
assign MEM[47714] = MEM[45561] + MEM[45616];
assign MEM[47715] = MEM[45562] + MEM[45641];
assign MEM[47716] = MEM[45563] + MEM[45617];
assign MEM[47717] = MEM[45564] + MEM[45606];
assign MEM[47718] = MEM[45565] + MEM[45590];
assign MEM[47719] = MEM[45571] + MEM[45743];
assign MEM[47720] = MEM[45573] + MEM[45636];
assign MEM[47721] = MEM[45578] + MEM[45649];
assign MEM[47722] = MEM[45579] + MEM[45669];
assign MEM[47723] = MEM[45581] + MEM[45646];
assign MEM[47724] = MEM[45582] + MEM[45638];
assign MEM[47725] = MEM[45583] + MEM[45621];
assign MEM[47726] = MEM[45585] + MEM[45607];
assign MEM[47727] = MEM[45586] + MEM[45595];
assign MEM[47728] = MEM[45587] + MEM[45618];
assign MEM[47729] = MEM[45591] + MEM[45655];
assign MEM[47730] = MEM[45592] + MEM[45630];
assign MEM[47731] = MEM[45593] + MEM[45687];
assign MEM[47732] = MEM[45596] + MEM[45662];
assign MEM[47733] = MEM[45598] + MEM[45639];
assign MEM[47734] = MEM[45599] + MEM[45626];
assign MEM[47735] = MEM[45600] + MEM[45719];
assign MEM[47736] = MEM[45601] + MEM[45654];
assign MEM[47737] = MEM[45602] + MEM[45678];
assign MEM[47738] = MEM[45609] + MEM[45685];
assign MEM[47739] = MEM[45611] + MEM[45660];
assign MEM[47740] = MEM[45612] + MEM[45632];
assign MEM[47741] = MEM[45619] + MEM[45675];
assign MEM[47742] = MEM[45622] + MEM[45691];
assign MEM[47743] = MEM[45623] + MEM[45762];
assign MEM[47744] = MEM[45624] + MEM[45724];
assign MEM[47745] = MEM[45625] + MEM[45701];
assign MEM[47746] = MEM[45628] + MEM[45652];
assign MEM[47747] = MEM[45629] + MEM[45707];
assign MEM[47748] = MEM[45631] + MEM[45792];
assign MEM[47749] = MEM[45634] + MEM[45684];
assign MEM[47750] = MEM[45635] + MEM[45704];
assign MEM[47751] = MEM[45637] + MEM[45674];
assign MEM[47752] = MEM[45640] + MEM[45759];
assign MEM[47753] = MEM[45642] + MEM[45712];
assign MEM[47754] = MEM[45643] + MEM[45700];
assign MEM[47755] = MEM[45644] + MEM[45695];
assign MEM[47756] = MEM[45645] + MEM[45754];
assign MEM[47757] = MEM[45648] + MEM[45698];
assign MEM[47758] = MEM[45650] + MEM[45697];
assign MEM[47759] = MEM[45651] + MEM[45716];
assign MEM[47760] = MEM[45653] + MEM[45677];
assign MEM[47761] = MEM[45656] + MEM[45689];
assign MEM[47762] = MEM[45657] + MEM[45705];
assign MEM[47763] = MEM[45658] + MEM[45692];
assign MEM[47764] = MEM[45659] + MEM[45746];
assign MEM[47765] = MEM[45661] + MEM[45738];
assign MEM[47766] = MEM[45664] + MEM[45690];
assign MEM[47767] = MEM[45666] + MEM[45715];
assign MEM[47768] = MEM[45667] + MEM[45773];
assign MEM[47769] = MEM[45668] + MEM[45725];
assign MEM[47770] = MEM[45670] + MEM[45713];
assign MEM[47771] = MEM[45671] + MEM[45777];
assign MEM[47772] = MEM[45672] + MEM[45751];
assign MEM[47773] = MEM[45676] + MEM[45745];
assign MEM[47774] = MEM[45679] + MEM[45714];
assign MEM[47775] = MEM[45680] + MEM[45750];
assign MEM[47776] = MEM[45681] + MEM[45729];
assign MEM[47777] = MEM[45682] + MEM[45744];
assign MEM[47778] = MEM[45683] + MEM[45748];
assign MEM[47779] = MEM[45686] + MEM[45717];
assign MEM[47780] = MEM[45688] + MEM[45736];
assign MEM[47781] = MEM[45693] + MEM[45735];
assign MEM[47782] = MEM[45694] + MEM[45742];
assign MEM[47783] = MEM[45699] + MEM[45732];
assign MEM[47784] = MEM[45702] + MEM[45793];
assign MEM[47785] = MEM[45703] + MEM[45741];
assign MEM[47786] = MEM[45706] + MEM[45780];
assign MEM[47787] = MEM[45708] + MEM[45730];
assign MEM[47788] = MEM[45709] + MEM[45737];
assign MEM[47789] = MEM[45710] + MEM[45782];
assign MEM[47790] = MEM[45711] + MEM[45761];
assign MEM[47791] = MEM[45718] + MEM[45813];
assign MEM[47792] = MEM[45720] + MEM[45826];
assign MEM[47793] = MEM[45721] + MEM[45784];
assign MEM[47794] = MEM[45722] + MEM[45829];
assign MEM[47795] = MEM[45723] + MEM[45837];
assign MEM[47796] = MEM[45726] + MEM[45766];
assign MEM[47797] = MEM[45727] + MEM[45756];
assign MEM[47798] = MEM[45728] + MEM[45814];
assign MEM[47799] = MEM[45731] + MEM[45786];
assign MEM[47800] = MEM[45733] + MEM[45802];
assign MEM[47801] = MEM[45734] + MEM[45875];
assign MEM[47802] = MEM[45739] + MEM[45767];
assign MEM[47803] = MEM[45740] + MEM[45816];
assign MEM[47804] = MEM[45747] + MEM[45874];
assign MEM[47805] = MEM[45749] + MEM[45817];
assign MEM[47806] = MEM[45752] + MEM[45809];
assign MEM[47807] = MEM[45753] + MEM[45785];
assign MEM[47808] = MEM[45755] + MEM[45808];
assign MEM[47809] = MEM[45757] + MEM[45800];
assign MEM[47810] = MEM[45758] + MEM[45889];
assign MEM[47811] = MEM[45760] + MEM[45805];
assign MEM[47812] = MEM[45763] + MEM[45783];
assign MEM[47813] = MEM[45764] + MEM[45798];
assign MEM[47814] = MEM[45765] + MEM[45840];
assign MEM[47815] = MEM[45768] + MEM[45852];
assign MEM[47816] = MEM[45769] + MEM[45797];
assign MEM[47817] = MEM[45770] + MEM[45832];
assign MEM[47818] = MEM[45771] + MEM[45833];
assign MEM[47819] = MEM[45772] + MEM[45855];
assign MEM[47820] = MEM[45774] + MEM[45863];
assign MEM[47821] = MEM[45775] + MEM[45861];
assign MEM[47822] = MEM[45776] + MEM[45827];
assign MEM[47823] = MEM[45778] + MEM[45828];
assign MEM[47824] = MEM[45779] + MEM[45881];
assign MEM[47825] = MEM[45781] + MEM[45865];
assign MEM[47826] = MEM[45787] + MEM[45853];
assign MEM[47827] = MEM[45788] + MEM[45838];
assign MEM[47828] = MEM[45789] + MEM[45845];
assign MEM[47829] = MEM[45790] + MEM[45841];
assign MEM[47830] = MEM[45791] + MEM[45880];
assign MEM[47831] = MEM[45794] + MEM[45892];
assign MEM[47832] = MEM[45795] + MEM[45862];
assign MEM[47833] = MEM[45796] + MEM[45896];
assign MEM[47834] = MEM[45799] + MEM[45834];
assign MEM[47835] = MEM[45801] + MEM[45859];
assign MEM[47836] = MEM[45803] + MEM[45847];
assign MEM[47837] = MEM[45804] + MEM[45849];
assign MEM[47838] = MEM[45806] + MEM[45903];
assign MEM[47839] = MEM[45807] + MEM[45836];
assign MEM[47840] = MEM[45810] + MEM[45906];
assign MEM[47841] = MEM[45811] + MEM[45877];
assign MEM[47842] = MEM[45812] + MEM[45885];
assign MEM[47843] = MEM[45815] + MEM[45898];
assign MEM[47844] = MEM[45818] + MEM[45842];
assign MEM[47845] = MEM[45819] + MEM[45868];
assign MEM[47846] = MEM[45820] + MEM[45844];
assign MEM[47847] = MEM[45821] + MEM[45856];
assign MEM[47848] = MEM[45822] + MEM[45894];
assign MEM[47849] = MEM[45823] + MEM[45860];
assign MEM[47850] = MEM[45824] + MEM[45895];
assign MEM[47851] = MEM[45825] + MEM[45901];
assign MEM[47852] = MEM[45830] + MEM[45883];
assign MEM[47853] = MEM[45831] + MEM[45893];
assign MEM[47854] = MEM[45835] + MEM[45887];
assign MEM[47855] = MEM[45839] + MEM[45907];
assign MEM[47856] = MEM[45843] + MEM[45940];
assign MEM[47857] = MEM[45846] + MEM[45870];
assign MEM[47858] = MEM[45848] + MEM[45912];
assign MEM[47859] = MEM[45850] + MEM[45932];
assign MEM[47860] = MEM[45851] + MEM[45867];
assign MEM[47861] = MEM[45854] + MEM[45899];
assign MEM[47862] = MEM[45857] + MEM[45948];
assign MEM[47863] = MEM[45858] + MEM[45917];
assign MEM[47864] = MEM[45864] + MEM[45965];
assign MEM[47865] = MEM[45866] + MEM[45905];
assign MEM[47866] = MEM[45869] + MEM[45956];
assign MEM[47867] = MEM[45871] + MEM[45934];
assign MEM[47868] = MEM[45872] + MEM[45921];
assign MEM[47869] = MEM[45873] + MEM[45949];
assign MEM[47870] = MEM[45876] + MEM[45961];
assign MEM[47871] = MEM[45878] + MEM[45967];
assign MEM[47872] = MEM[45879] + MEM[45922];
assign MEM[47873] = MEM[45882] + MEM[45909];
assign MEM[47874] = MEM[45884] + MEM[45947];
assign MEM[47875] = MEM[45886] + MEM[45958];
assign MEM[47876] = MEM[45888] + MEM[45980];
assign MEM[47877] = MEM[45890] + MEM[45976];
assign MEM[47878] = MEM[45891] + MEM[45944];
assign MEM[47879] = MEM[45897] + MEM[45927];
assign MEM[47880] = MEM[45900] + MEM[45928];
assign MEM[47881] = MEM[45902] + MEM[45986];
assign MEM[47882] = MEM[45904] + MEM[45974];
assign MEM[47883] = MEM[45908] + MEM[45988];
assign MEM[47884] = MEM[45910] + MEM[45972];
assign MEM[47885] = MEM[45911] + MEM[45966];
assign MEM[47886] = MEM[45913] + MEM[45992];
assign MEM[47887] = MEM[45914] + MEM[45981];
assign MEM[47888] = MEM[45915] + MEM[46044];
assign MEM[47889] = MEM[45916] + MEM[46004];
assign MEM[47890] = MEM[45918] + MEM[45993];
assign MEM[47891] = MEM[45919] + MEM[46013];
assign MEM[47892] = MEM[45920] + MEM[46008];
assign MEM[47893] = MEM[45923] + MEM[46000];
assign MEM[47894] = MEM[45924] + MEM[46039];
assign MEM[47895] = MEM[45925] + MEM[45982];
assign MEM[47896] = MEM[45926] + MEM[45994];
assign MEM[47897] = MEM[45929] + MEM[45983];
assign MEM[47898] = MEM[45930] + MEM[45943];
assign MEM[47899] = MEM[45931] + MEM[46050];
assign MEM[47900] = MEM[45933] + MEM[45954];
assign MEM[47901] = MEM[45935] + MEM[45971];
assign MEM[47902] = MEM[45936] + MEM[45984];
assign MEM[47903] = MEM[45937] + MEM[46005];
assign MEM[47904] = MEM[45938] + MEM[45990];
assign MEM[47905] = MEM[45939] + MEM[46031];
assign MEM[47906] = MEM[45941] + MEM[45991];
assign MEM[47907] = MEM[45942] + MEM[45998];
assign MEM[47908] = MEM[45945] + MEM[45999];
assign MEM[47909] = MEM[45946] + MEM[45979];
assign MEM[47910] = MEM[45950] + MEM[46018];
assign MEM[47911] = MEM[45951] + MEM[46106];
assign MEM[47912] = MEM[45952] + MEM[46002];
assign MEM[47913] = MEM[45953] + MEM[46006];
assign MEM[47914] = MEM[45955] + MEM[46025];
assign MEM[47915] = MEM[45957] + MEM[46024];
assign MEM[47916] = MEM[45959] + MEM[45987];
assign MEM[47917] = MEM[45960] + MEM[46011];
assign MEM[47918] = MEM[45962] + MEM[45975];
assign MEM[47919] = MEM[45963] + MEM[46014];
assign MEM[47920] = MEM[45964] + MEM[46027];
assign MEM[47921] = MEM[45968] + MEM[46003];
assign MEM[47922] = MEM[45969] + MEM[46043];
assign MEM[47923] = MEM[45970] + MEM[45997];
assign MEM[47924] = MEM[45973] + MEM[46007];
assign MEM[47925] = MEM[45977] + MEM[46019];
assign MEM[47926] = MEM[45978] + MEM[46026];
assign MEM[47927] = MEM[45985] + MEM[46072];
assign MEM[47928] = MEM[45989] + MEM[46073];
assign MEM[47929] = MEM[45995] + MEM[46030];
assign MEM[47930] = MEM[45996] + MEM[46089];
assign MEM[47931] = MEM[46001] + MEM[46075];
assign MEM[47932] = MEM[46009] + MEM[46058];
assign MEM[47933] = MEM[46010] + MEM[46076];
assign MEM[47934] = MEM[46012] + MEM[46081];
assign MEM[47935] = MEM[46015] + MEM[46086];
assign MEM[47936] = MEM[46016] + MEM[46082];
assign MEM[47937] = MEM[46017] + MEM[46057];
assign MEM[47938] = MEM[46020] + MEM[46036];
assign MEM[47939] = MEM[46021] + MEM[46097];
assign MEM[47940] = MEM[46022] + MEM[46077];
assign MEM[47941] = MEM[46023] + MEM[46122];
assign MEM[47942] = MEM[46028] + MEM[46110];
assign MEM[47943] = MEM[46029] + MEM[46078];
assign MEM[47944] = MEM[46032] + MEM[46189];
assign MEM[47945] = MEM[46033] + MEM[46116];
assign MEM[47946] = MEM[46034] + MEM[46108];
assign MEM[47947] = MEM[46035] + MEM[46079];
assign MEM[47948] = MEM[46037] + MEM[46099];
assign MEM[47949] = MEM[46038] + MEM[46114];
assign MEM[47950] = MEM[46040] + MEM[46095];
assign MEM[47951] = MEM[46041] + MEM[46094];
assign MEM[47952] = MEM[46042] + MEM[46098];
assign MEM[47953] = MEM[46045] + MEM[46069];
assign MEM[47954] = MEM[46046] + MEM[46123];
assign MEM[47955] = MEM[46047] + MEM[46133];
assign MEM[47956] = MEM[46048] + MEM[46136];
assign MEM[47957] = MEM[46049] + MEM[46084];
assign MEM[47958] = MEM[46051] + MEM[46091];
assign MEM[47959] = MEM[46052] + MEM[46103];
assign MEM[47960] = MEM[46053] + MEM[46104];
assign MEM[47961] = MEM[46054] + MEM[46090];
assign MEM[47962] = MEM[46055] + MEM[46170];
assign MEM[47963] = MEM[46056] + MEM[46128];
assign MEM[47964] = MEM[46059] + MEM[46144];
assign MEM[47965] = MEM[46060] + MEM[46125];
assign MEM[47966] = MEM[46061] + MEM[46142];
assign MEM[47967] = MEM[46062] + MEM[46134];
assign MEM[47968] = MEM[46063] + MEM[46141];
assign MEM[47969] = MEM[46064] + MEM[46109];
assign MEM[47970] = MEM[46065] + MEM[46143];
assign MEM[47971] = MEM[46066] + MEM[46139];
assign MEM[47972] = MEM[46067] + MEM[46188];
assign MEM[47973] = MEM[46068] + MEM[46124];
assign MEM[47974] = MEM[46070] + MEM[46127];
assign MEM[47975] = MEM[46071] + MEM[46149];
assign MEM[47976] = MEM[46074] + MEM[46150];
assign MEM[47977] = MEM[46080] + MEM[46151];
assign MEM[47978] = MEM[46083] + MEM[46183];
assign MEM[47979] = MEM[46085] + MEM[46138];
assign MEM[47980] = MEM[46087] + MEM[46115];
assign MEM[47981] = MEM[46088] + MEM[46165];
assign MEM[47982] = MEM[46092] + MEM[46154];
assign MEM[47983] = MEM[46093] + MEM[46163];
assign MEM[47984] = MEM[46096] + MEM[46156];
assign MEM[47985] = MEM[46100] + MEM[46177];
assign MEM[47986] = MEM[46101] + MEM[46146];
assign MEM[47987] = MEM[46102] + MEM[46179];
assign MEM[47988] = MEM[46105] + MEM[46157];
assign MEM[47989] = MEM[46107] + MEM[46187];
assign MEM[47990] = MEM[46111] + MEM[46198];
assign MEM[47991] = MEM[46112] + MEM[46186];
assign MEM[47992] = MEM[46113] + MEM[46180];
assign MEM[47993] = MEM[46117] + MEM[46168];
assign MEM[47994] = MEM[46118] + MEM[46226];
assign MEM[47995] = MEM[46119] + MEM[46199];
assign MEM[47996] = MEM[46120] + MEM[46206];
assign MEM[47997] = MEM[46121] + MEM[46178];
assign MEM[47998] = MEM[46126] + MEM[46223];
assign MEM[47999] = MEM[46129] + MEM[46209];
assign MEM[48000] = MEM[46130] + MEM[46182];
assign MEM[48001] = MEM[46131] + MEM[46197];
assign MEM[48002] = MEM[46132] + MEM[46241];
assign MEM[48003] = MEM[46135] + MEM[46175];
assign MEM[48004] = MEM[46137] + MEM[46176];
assign MEM[48005] = MEM[46140] + MEM[46210];
assign MEM[48006] = MEM[46145] + MEM[46255];
assign MEM[48007] = MEM[46147] + MEM[46219];
assign MEM[48008] = MEM[46148] + MEM[46248];
assign MEM[48009] = MEM[46152] + MEM[46216];
assign MEM[48010] = MEM[46153] + MEM[46194];
assign MEM[48011] = MEM[46155] + MEM[46244];
assign MEM[48012] = MEM[46158] + MEM[46203];
assign MEM[48013] = MEM[46159] + MEM[46218];
assign MEM[48014] = MEM[46160] + MEM[46201];
assign MEM[48015] = MEM[46161] + MEM[46232];
assign MEM[48016] = MEM[46162] + MEM[46192];
assign MEM[48017] = MEM[46164] + MEM[46266];
assign MEM[48018] = MEM[46166] + MEM[46208];
assign MEM[48019] = MEM[46167] + MEM[46222];
assign MEM[48020] = MEM[46169] + MEM[46234];
assign MEM[48021] = MEM[46171] + MEM[46221];
assign MEM[48022] = MEM[46172] + MEM[46227];
assign MEM[48023] = MEM[46173] + MEM[46238];
assign MEM[48024] = MEM[46174] + MEM[46207];
assign MEM[48025] = MEM[46181] + MEM[46233];
assign MEM[48026] = MEM[46184] + MEM[46225];
assign MEM[48027] = MEM[46185] + MEM[46217];
assign MEM[48028] = MEM[46190] + MEM[46269];
assign MEM[48029] = MEM[46191] + MEM[46242];
assign MEM[48030] = MEM[46193] + MEM[46259];
assign MEM[48031] = MEM[46195] + MEM[46247];
assign MEM[48032] = MEM[46196] + MEM[46271];
assign MEM[48033] = MEM[46200] + MEM[46254];
assign MEM[48034] = MEM[46202] + MEM[46264];
assign MEM[48035] = MEM[46204] + MEM[46246];
assign MEM[48036] = MEM[46205] + MEM[46257];
assign MEM[48037] = MEM[46211] + MEM[46272];
assign MEM[48038] = MEM[46212] + MEM[46270];
assign MEM[48039] = MEM[46213] + MEM[46260];
assign MEM[48040] = MEM[46214] + MEM[46306];
assign MEM[48041] = MEM[46215] + MEM[46277];
assign MEM[48042] = MEM[46220] + MEM[46279];
assign MEM[48043] = MEM[46224] + MEM[46313];
assign MEM[48044] = MEM[46228] + MEM[46295];
assign MEM[48045] = MEM[46229] + MEM[46315];
assign MEM[48046] = MEM[46230] + MEM[46263];
assign MEM[48047] = MEM[46231] + MEM[46339];
assign MEM[48048] = MEM[46235] + MEM[46314];
assign MEM[48049] = MEM[46236] + MEM[46329];
assign MEM[48050] = MEM[46237] + MEM[46293];
assign MEM[48051] = MEM[46239] + MEM[46334];
assign MEM[48052] = MEM[46240] + MEM[46298];
assign MEM[48053] = MEM[46243] + MEM[46325];
assign MEM[48054] = MEM[46245] + MEM[46288];
assign MEM[48055] = MEM[46249] + MEM[46341];
assign MEM[48056] = MEM[46250] + MEM[46283];
assign MEM[48057] = MEM[46251] + MEM[46285];
assign MEM[48058] = MEM[46252] + MEM[46395];
assign MEM[48059] = MEM[46253] + MEM[46300];
assign MEM[48060] = MEM[46256] + MEM[46303];
assign MEM[48061] = MEM[46258] + MEM[46311];
assign MEM[48062] = MEM[46261] + MEM[46324];
assign MEM[48063] = MEM[46262] + MEM[46321];
assign MEM[48064] = MEM[46265] + MEM[46331];
assign MEM[48065] = MEM[46267] + MEM[46364];
assign MEM[48066] = MEM[46268] + MEM[46317];
assign MEM[48067] = MEM[46273] + MEM[46345];
assign MEM[48068] = MEM[46274] + MEM[46319];
assign MEM[48069] = MEM[46275] + MEM[46342];
assign MEM[48070] = MEM[46276] + MEM[46337];
assign MEM[48071] = MEM[46278] + MEM[46336];
assign MEM[48072] = MEM[46280] + MEM[46379];
assign MEM[48073] = MEM[46281] + MEM[46389];
assign MEM[48074] = MEM[46282] + MEM[46310];
assign MEM[48075] = MEM[46284] + MEM[46340];
assign MEM[48076] = MEM[46286] + MEM[46349];
assign MEM[48077] = MEM[46287] + MEM[46347];
assign MEM[48078] = MEM[46289] + MEM[46350];
assign MEM[48079] = MEM[46290] + MEM[46352];
assign MEM[48080] = MEM[46291] + MEM[46377];
assign MEM[48081] = MEM[46292] + MEM[46338];
assign MEM[48082] = MEM[46294] + MEM[46380];
assign MEM[48083] = MEM[46296] + MEM[46326];
assign MEM[48084] = MEM[46297] + MEM[46398];
assign MEM[48085] = MEM[46299] + MEM[46406];
assign MEM[48086] = MEM[46301] + MEM[46343];
assign MEM[48087] = MEM[46302] + MEM[46358];
assign MEM[48088] = MEM[46304] + MEM[46371];
assign MEM[48089] = MEM[46305] + MEM[46366];
assign MEM[48090] = MEM[46307] + MEM[46346];
assign MEM[48091] = MEM[46308] + MEM[46399];
assign MEM[48092] = MEM[46309] + MEM[46363];
assign MEM[48093] = MEM[46312] + MEM[46375];
assign MEM[48094] = MEM[46316] + MEM[46359];
assign MEM[48095] = MEM[46318] + MEM[46477];
assign MEM[48096] = MEM[46320] + MEM[46423];
assign MEM[48097] = MEM[46322] + MEM[46370];
assign MEM[48098] = MEM[46323] + MEM[46382];
assign MEM[48099] = MEM[46327] + MEM[46392];
assign MEM[48100] = MEM[46328] + MEM[46361];
assign MEM[48101] = MEM[46330] + MEM[46372];
assign MEM[48102] = MEM[46332] + MEM[46425];
assign MEM[48103] = MEM[46333] + MEM[46368];
assign MEM[48104] = MEM[46335] + MEM[46402];
assign MEM[48105] = MEM[46344] + MEM[46426];
assign MEM[48106] = MEM[46348] + MEM[46384];
assign MEM[48107] = MEM[46351] + MEM[46415];
assign MEM[48108] = MEM[46353] + MEM[46411];
assign MEM[48109] = MEM[46354] + MEM[46438];
assign MEM[48110] = MEM[46355] + MEM[46397];
assign MEM[48111] = MEM[46356] + MEM[46409];
assign MEM[48112] = MEM[46357] + MEM[46432];
assign MEM[48113] = MEM[46360] + MEM[46422];
assign MEM[48114] = MEM[46362] + MEM[46437];
assign MEM[48115] = MEM[46365] + MEM[46435];
assign MEM[48116] = MEM[46367] + MEM[46421];
assign MEM[48117] = MEM[46369] + MEM[46453];
assign MEM[48118] = MEM[46373] + MEM[46478];
assign MEM[48119] = MEM[46374] + MEM[46441];
assign MEM[48120] = MEM[46376] + MEM[46483];
assign MEM[48121] = MEM[46378] + MEM[46427];
assign MEM[48122] = MEM[46381] + MEM[46462];
assign MEM[48123] = MEM[46383] + MEM[46442];
assign MEM[48124] = MEM[46385] + MEM[46451];
assign MEM[48125] = MEM[46386] + MEM[46443];
assign MEM[48126] = MEM[46387] + MEM[46463];
assign MEM[48127] = MEM[46388] + MEM[46431];
assign MEM[48128] = MEM[46390] + MEM[46450];
assign MEM[48129] = MEM[46391] + MEM[46448];
assign MEM[48130] = MEM[46393] + MEM[46459];
assign MEM[48131] = MEM[46394] + MEM[46455];
assign MEM[48132] = MEM[46396] + MEM[46454];
assign MEM[48133] = MEM[46400] + MEM[46428];
assign MEM[48134] = MEM[46401] + MEM[46473];
assign MEM[48135] = MEM[46403] + MEM[46467];
assign MEM[48136] = MEM[46404] + MEM[46444];
assign MEM[48137] = MEM[46405] + MEM[46457];
assign MEM[48138] = MEM[46407] + MEM[46468];
assign MEM[48139] = MEM[46408] + MEM[46445];
assign MEM[48140] = MEM[46410] + MEM[46475];
assign MEM[48141] = MEM[46412] + MEM[46505];
assign MEM[48142] = MEM[46413] + MEM[46436];
assign MEM[48143] = MEM[46414] + MEM[46479];
assign MEM[48144] = MEM[46416] + MEM[46508];
assign MEM[48145] = MEM[46417] + MEM[46492];
assign MEM[48146] = MEM[46418] + MEM[46460];
assign MEM[48147] = MEM[46419] + MEM[46476];
assign MEM[48148] = MEM[46420] + MEM[46474];
assign MEM[48149] = MEM[46424] + MEM[46499];
assign MEM[48150] = MEM[46429] + MEM[46494];
assign MEM[48151] = MEM[46430] + MEM[46514];
assign MEM[48152] = MEM[46433] + MEM[46512];
assign MEM[48153] = MEM[46434] + MEM[46484];
assign MEM[48154] = MEM[46439] + MEM[46510];
assign MEM[48155] = MEM[46440] + MEM[46509];
assign MEM[48156] = MEM[46446] + MEM[46471];
assign MEM[48157] = MEM[46447] + MEM[46500];
assign MEM[48158] = MEM[46449] + MEM[46527];
assign MEM[48159] = MEM[46452] + MEM[46529];
assign MEM[48160] = MEM[46456] + MEM[46525];
assign MEM[48161] = MEM[46458] + MEM[46504];
assign MEM[48162] = MEM[46461] + MEM[46542];
assign MEM[48163] = MEM[46464] + MEM[46534];
assign MEM[48164] = MEM[46465] + MEM[46531];
assign MEM[48165] = MEM[46466] + MEM[46536];
assign MEM[48166] = MEM[46469] + MEM[46507];
assign MEM[48167] = MEM[46470] + MEM[46498];
assign MEM[48168] = MEM[46472] + MEM[46511];
assign MEM[48169] = MEM[46480] + MEM[46550];
assign MEM[48170] = MEM[46481] + MEM[46543];
assign MEM[48171] = MEM[46482] + MEM[46547];
assign MEM[48172] = MEM[46485] + MEM[46532];
assign MEM[48173] = MEM[46486] + MEM[46579];
assign MEM[48174] = MEM[46487] + MEM[46557];
assign MEM[48175] = MEM[46488] + MEM[46574];
assign MEM[48176] = MEM[46489] + MEM[46558];
assign MEM[48177] = MEM[46490] + MEM[46544];
assign MEM[48178] = MEM[46491] + MEM[46539];
assign MEM[48179] = MEM[46493] + MEM[46548];
assign MEM[48180] = MEM[46495] + MEM[46566];
assign MEM[48181] = MEM[46496] + MEM[46564];
assign MEM[48182] = MEM[46497] + MEM[46535];
assign MEM[48183] = MEM[46501] + MEM[46584];
assign MEM[48184] = MEM[46502] + MEM[46618];
assign MEM[48185] = MEM[46503] + MEM[46538];
assign MEM[48186] = MEM[46506] + MEM[46545];
assign MEM[48187] = MEM[46513] + MEM[46552];
assign MEM[48188] = MEM[46515] + MEM[46591];
assign MEM[48189] = MEM[46516] + MEM[46571];
assign MEM[48190] = MEM[46517] + MEM[46616];
assign MEM[48191] = MEM[46518] + MEM[46657];
assign MEM[48192] = MEM[46519] + MEM[46643];
assign MEM[48193] = MEM[46520] + MEM[46581];
assign MEM[48194] = MEM[46521] + MEM[46597];
assign MEM[48195] = MEM[46522] + MEM[46596];
assign MEM[48196] = MEM[46523] + MEM[46572];
assign MEM[48197] = MEM[46524] + MEM[46576];
assign MEM[48198] = MEM[46526] + MEM[46561];
assign MEM[48199] = MEM[46528] + MEM[46575];
assign MEM[48200] = MEM[46530] + MEM[46582];
assign MEM[48201] = MEM[46533] + MEM[46563];
assign MEM[48202] = MEM[46537] + MEM[46570];
assign MEM[48203] = MEM[46540] + MEM[46588];
assign MEM[48204] = MEM[46541] + MEM[46567];
assign MEM[48205] = MEM[46546] + MEM[46603];
assign MEM[48206] = MEM[46549] + MEM[46628];
assign MEM[48207] = MEM[46551] + MEM[46583];
assign MEM[48208] = MEM[46553] + MEM[46636];
assign MEM[48209] = MEM[46554] + MEM[46605];
assign MEM[48210] = MEM[46555] + MEM[46610];
assign MEM[48211] = MEM[46556] + MEM[46595];
assign MEM[48212] = MEM[46559] + MEM[46633];
assign MEM[48213] = MEM[46560] + MEM[46606];
assign MEM[48214] = MEM[46562] + MEM[46609];
assign MEM[48215] = MEM[46565] + MEM[46667];
assign MEM[48216] = MEM[46568] + MEM[46625];
assign MEM[48217] = MEM[46569] + MEM[46614];
assign MEM[48218] = MEM[46573] + MEM[46611];
assign MEM[48219] = MEM[46577] + MEM[46602];
assign MEM[48220] = MEM[46578] + MEM[46634];
assign MEM[48221] = MEM[46580] + MEM[46644];
assign MEM[48222] = MEM[46585] + MEM[46632];
assign MEM[48223] = MEM[46586] + MEM[46630];
assign MEM[48224] = MEM[46587] + MEM[46672];
assign MEM[48225] = MEM[46589] + MEM[46629];
assign MEM[48226] = MEM[46590] + MEM[46647];
assign MEM[48227] = MEM[46592] + MEM[46640];
assign MEM[48228] = MEM[46593] + MEM[46658];
assign MEM[48229] = MEM[46594] + MEM[46665];
assign MEM[48230] = MEM[46598] + MEM[46661];
assign MEM[48231] = MEM[46599] + MEM[46678];
assign MEM[48232] = MEM[46600] + MEM[46656];
assign MEM[48233] = MEM[46601] + MEM[46682];
assign MEM[48234] = MEM[46604] + MEM[46655];
assign MEM[48235] = MEM[46607] + MEM[46666];
assign MEM[48236] = MEM[46608] + MEM[46675];
assign MEM[48237] = MEM[46612] + MEM[46684];
assign MEM[48238] = MEM[46613] + MEM[46652];
assign MEM[48239] = MEM[46615] + MEM[46668];
assign MEM[48240] = MEM[46617] + MEM[46720];
assign MEM[48241] = MEM[46619] + MEM[46714];
assign MEM[48242] = MEM[46620] + MEM[46685];
assign MEM[48243] = MEM[46621] + MEM[46749];
assign MEM[48244] = MEM[46622] + MEM[46681];
assign MEM[48245] = MEM[46623] + MEM[46687];
assign MEM[48246] = MEM[46624] + MEM[46700];
assign MEM[48247] = MEM[46626] + MEM[46669];
assign MEM[48248] = MEM[46627] + MEM[46688];
assign MEM[48249] = MEM[46631] + MEM[46702];
assign MEM[48250] = MEM[46635] + MEM[46680];
assign MEM[48251] = MEM[46637] + MEM[46677];
assign MEM[48252] = MEM[46638] + MEM[46683];
assign MEM[48253] = MEM[46639] + MEM[46716];
assign MEM[48254] = MEM[46641] + MEM[46691];
assign MEM[48255] = MEM[46642] + MEM[46701];
assign MEM[48256] = MEM[46645] + MEM[46696];
assign MEM[48257] = MEM[46646] + MEM[46738];
assign MEM[48258] = MEM[46648] + MEM[46731];
assign MEM[48259] = MEM[46649] + MEM[46763];
assign MEM[48260] = MEM[46650] + MEM[46722];
assign MEM[48261] = MEM[46651] + MEM[46709];
assign MEM[48262] = MEM[46653] + MEM[46694];
assign MEM[48263] = MEM[46654] + MEM[46697];
assign MEM[48264] = MEM[46659] + MEM[46726];
assign MEM[48265] = MEM[46660] + MEM[46721];
assign MEM[48266] = MEM[46662] + MEM[46689];
assign MEM[48267] = MEM[46663] + MEM[46718];
assign MEM[48268] = MEM[46664] + MEM[46737];
assign MEM[48269] = MEM[46670] + MEM[46740];
assign MEM[48270] = MEM[46671] + MEM[46748];
assign MEM[48271] = MEM[46673] + MEM[46733];
assign MEM[48272] = MEM[46674] + MEM[46686];
assign MEM[48273] = MEM[46676] + MEM[46710];
assign MEM[48274] = MEM[46679] + MEM[46766];
assign MEM[48275] = MEM[46690] + MEM[46727];
assign MEM[48276] = MEM[46692] + MEM[46769];
assign MEM[48277] = MEM[46693] + MEM[46779];
assign MEM[48278] = MEM[46695] + MEM[46790];
assign MEM[48279] = MEM[46698] + MEM[46780];
assign MEM[48280] = MEM[46699] + MEM[46764];
assign MEM[48281] = MEM[46703] + MEM[46776];
assign MEM[48282] = MEM[46704] + MEM[46746];
assign MEM[48283] = MEM[46705] + MEM[46768];
assign MEM[48284] = MEM[46706] + MEM[46810];
assign MEM[48285] = MEM[46707] + MEM[46755];
assign MEM[48286] = MEM[46708] + MEM[46774];
assign MEM[48287] = MEM[46711] + MEM[46775];
assign MEM[48288] = MEM[46712] + MEM[46814];
assign MEM[48289] = MEM[46713] + MEM[46778];
assign MEM[48290] = MEM[46715] + MEM[46786];
assign MEM[48291] = MEM[46717] + MEM[46794];
assign MEM[48292] = MEM[46719] + MEM[46758];
assign MEM[48293] = MEM[46723] + MEM[46813];
assign MEM[48294] = MEM[46724] + MEM[46804];
assign MEM[48295] = MEM[46725] + MEM[46805];
assign MEM[48296] = MEM[46728] + MEM[46793];
assign MEM[48297] = MEM[46729] + MEM[46807];
assign MEM[48298] = MEM[46730] + MEM[46773];
assign MEM[48299] = MEM[46732] + MEM[46815];
assign MEM[48300] = MEM[46734] + MEM[46820];
assign MEM[48301] = MEM[46735] + MEM[46785];
assign MEM[48302] = MEM[46736] + MEM[46762];
assign MEM[48303] = MEM[46739] + MEM[46825];
assign MEM[48304] = MEM[46741] + MEM[46782];
assign MEM[48305] = MEM[46742] + MEM[46818];
assign MEM[48306] = MEM[46743] + MEM[46827];
assign MEM[48307] = MEM[46744] + MEM[46802];
assign MEM[48308] = MEM[46745] + MEM[46795];
assign MEM[48309] = MEM[46747] + MEM[46777];
assign MEM[48310] = MEM[46750] + MEM[46781];
assign MEM[48311] = MEM[46751] + MEM[46792];
assign MEM[48312] = MEM[46752] + MEM[46809];
assign MEM[48313] = MEM[46753] + MEM[46840];
assign MEM[48314] = MEM[46754] + MEM[46828];
assign MEM[48315] = MEM[46756] + MEM[46812];
assign MEM[48316] = MEM[46757] + MEM[46858];
assign MEM[48317] = MEM[46759] + MEM[46801];
assign MEM[48318] = MEM[46760] + MEM[46799];
assign MEM[48319] = MEM[46761] + MEM[46834];
assign MEM[48320] = MEM[46765] + MEM[46845];
assign MEM[48321] = MEM[46767] + MEM[46843];
assign MEM[48322] = MEM[46770] + MEM[46808];
assign MEM[48323] = MEM[46771] + MEM[46839];
assign MEM[48324] = MEM[46772] + MEM[46849];
assign MEM[48325] = MEM[46783] + MEM[46841];
assign MEM[48326] = MEM[46784] + MEM[46874];
assign MEM[48327] = MEM[46787] + MEM[46867];
assign MEM[48328] = MEM[46788] + MEM[46824];
assign MEM[48329] = MEM[46789] + MEM[46835];
assign MEM[48330] = MEM[46791] + MEM[46879];
assign MEM[48331] = MEM[46796] + MEM[46844];
assign MEM[48332] = MEM[46797] + MEM[46926];
assign MEM[48333] = MEM[46798] + MEM[46881];
assign MEM[48334] = MEM[46800] + MEM[46880];
assign MEM[48335] = MEM[46803] + MEM[46887];
assign MEM[48336] = MEM[46806] + MEM[46866];
assign MEM[48337] = MEM[46811] + MEM[46853];
assign MEM[48338] = MEM[46816] + MEM[46863];
assign MEM[48339] = MEM[46817] + MEM[46847];
assign MEM[48340] = MEM[46819] + MEM[46861];
assign MEM[48341] = MEM[46821] + MEM[46872];
assign MEM[48342] = MEM[46822] + MEM[46891];
assign MEM[48343] = MEM[46823] + MEM[46873];
assign MEM[48344] = MEM[46826] + MEM[46959];
assign MEM[48345] = MEM[46829] + MEM[46868];
assign MEM[48346] = MEM[46830] + MEM[46893];
assign MEM[48347] = MEM[46831] + MEM[46912];
assign MEM[48348] = MEM[46832] + MEM[46877];
assign MEM[48349] = MEM[46833] + MEM[46901];
assign MEM[48350] = MEM[46836] + MEM[46932];
assign MEM[48351] = MEM[46837] + MEM[46876];
assign MEM[48352] = MEM[46838] + MEM[46914];
assign MEM[48353] = MEM[46842] + MEM[46902];
assign MEM[48354] = MEM[46846] + MEM[46870];
assign MEM[48355] = MEM[46848] + MEM[46903];
assign MEM[48356] = MEM[46850] + MEM[46897];
assign MEM[48357] = MEM[46851] + MEM[46931];
assign MEM[48358] = MEM[46852] + MEM[46915];
assign MEM[48359] = MEM[46854] + MEM[46922];
assign MEM[48360] = MEM[46855] + MEM[46957];
assign MEM[48361] = MEM[46856] + MEM[46930];
assign MEM[48362] = MEM[46857] + MEM[46898];
assign MEM[48363] = MEM[46859] + MEM[46904];
assign MEM[48364] = MEM[46860] + MEM[46910];
assign MEM[48365] = MEM[46862] + MEM[46900];
assign MEM[48366] = MEM[46864] + MEM[46896];
assign MEM[48367] = MEM[46865] + MEM[46974];
assign MEM[48368] = MEM[46869] + MEM[46940];
assign MEM[48369] = MEM[46871] + MEM[46923];
assign MEM[48370] = MEM[46875] + MEM[46935];
assign MEM[48371] = MEM[46878] + MEM[46929];
assign MEM[48372] = MEM[46882] + MEM[46920];
assign MEM[48373] = MEM[46883] + MEM[46945];
assign MEM[48374] = MEM[46884] + MEM[46970];
assign MEM[48375] = MEM[46885] + MEM[46938];
assign MEM[48376] = MEM[46886] + MEM[46956];
assign MEM[48377] = MEM[46888] + MEM[46961];
assign MEM[48378] = MEM[46889] + MEM[46925];
assign MEM[48379] = MEM[46890] + MEM[46949];
assign MEM[48380] = MEM[46892] + MEM[46976];
assign MEM[48381] = MEM[46894] + MEM[46917];
assign MEM[48382] = MEM[46895] + MEM[46972];
assign MEM[48383] = MEM[46899] + MEM[46947];
assign MEM[48384] = MEM[46905] + MEM[47017];
assign MEM[48385] = MEM[46906] + MEM[46962];
assign MEM[48386] = MEM[46907] + MEM[46975];
assign MEM[48387] = MEM[46908] + MEM[46971];
assign MEM[48388] = MEM[46909] + MEM[46969];
assign MEM[48389] = MEM[46911] + MEM[46953];
assign MEM[48390] = MEM[46913] + MEM[46952];
assign MEM[48391] = MEM[46916] + MEM[46984];
assign MEM[48392] = MEM[46918] + MEM[46937];
assign MEM[48393] = MEM[46919] + MEM[46980];
assign MEM[48394] = MEM[46921] + MEM[47002];
assign MEM[48395] = MEM[46924] + MEM[46994];
assign MEM[48396] = MEM[46927] + MEM[47015];
assign MEM[48397] = MEM[46928] + MEM[47022];
assign MEM[48398] = MEM[46933] + MEM[46991];
assign MEM[48399] = MEM[46934] + MEM[46966];
assign MEM[48400] = MEM[46936] + MEM[46996];
assign MEM[48401] = MEM[46939] + MEM[46987];
assign MEM[48402] = MEM[46941] + MEM[46988];
assign MEM[48403] = MEM[46942] + MEM[47006];
assign MEM[48404] = MEM[46943] + MEM[47011];
assign MEM[48405] = MEM[46944] + MEM[47013];
assign MEM[48406] = MEM[46946] + MEM[47010];
assign MEM[48407] = MEM[46948] + MEM[47028];
assign MEM[48408] = MEM[46950] + MEM[47020];
assign MEM[48409] = MEM[46951] + MEM[46982];
assign MEM[48410] = MEM[46954] + MEM[47019];
assign MEM[48411] = MEM[46955] + MEM[47005];
assign MEM[48412] = MEM[46958] + MEM[47004];
assign MEM[48413] = MEM[46960] + MEM[47014];
assign MEM[48414] = MEM[46963] + MEM[47026];
assign MEM[48415] = MEM[46964] + MEM[47068];
assign MEM[48416] = MEM[46965] + MEM[47040];
assign MEM[48417] = MEM[46967] + MEM[47001];
assign MEM[48418] = MEM[46968] + MEM[47076];
assign MEM[48419] = MEM[46973] + MEM[47037];
assign MEM[48420] = MEM[46977] + MEM[47072];
assign MEM[48421] = MEM[46978] + MEM[47033];
assign MEM[48422] = MEM[46979] + MEM[47025];
assign MEM[48423] = MEM[46981] + MEM[47049];
assign MEM[48424] = MEM[46983] + MEM[47066];
assign MEM[48425] = MEM[46985] + MEM[47048];
assign MEM[48426] = MEM[46986] + MEM[47043];
assign MEM[48427] = MEM[46989] + MEM[47035];
assign MEM[48428] = MEM[46990] + MEM[47007];
assign MEM[48429] = MEM[46992] + MEM[47050];
assign MEM[48430] = MEM[46993] + MEM[47041];
assign MEM[48431] = MEM[46995] + MEM[47082];
assign MEM[48432] = MEM[46997] + MEM[47051];
assign MEM[48433] = MEM[46998] + MEM[47052];
assign MEM[48434] = MEM[46999] + MEM[47047];
assign MEM[48435] = MEM[47000] + MEM[47055];
assign MEM[48436] = MEM[47003] + MEM[47081];
assign MEM[48437] = MEM[47008] + MEM[47044];
assign MEM[48438] = MEM[47009] + MEM[47065];
assign MEM[48439] = MEM[47012] + MEM[47092];
assign MEM[48440] = MEM[47016] + MEM[47079];
assign MEM[48441] = MEM[47018] + MEM[47083];
assign MEM[48442] = MEM[47021] + MEM[47078];
assign MEM[48443] = MEM[47023] + MEM[47088];
assign MEM[48444] = MEM[47024] + MEM[47125];
assign MEM[48445] = MEM[47027] + MEM[47102];
assign MEM[48446] = MEM[47029] + MEM[47107];
assign MEM[48447] = MEM[47030] + MEM[47115];
assign MEM[48448] = MEM[47031] + MEM[47108];
assign MEM[48449] = MEM[47032] + MEM[47109];
assign MEM[48450] = MEM[47034] + MEM[47090];
assign MEM[48451] = MEM[47036] + MEM[47126];
assign MEM[48452] = MEM[47038] + MEM[47111];
assign MEM[48453] = MEM[47039] + MEM[47086];
assign MEM[48454] = MEM[47042] + MEM[47073];
assign MEM[48455] = MEM[47045] + MEM[47121];
assign MEM[48456] = MEM[47046] + MEM[47144];
assign MEM[48457] = MEM[47053] + MEM[47127];
assign MEM[48458] = MEM[47054] + MEM[47106];
assign MEM[48459] = MEM[47056] + MEM[47100];
assign MEM[48460] = MEM[47057] + MEM[47148];
assign MEM[48461] = MEM[47058] + MEM[47129];
assign MEM[48462] = MEM[47059] + MEM[47114];
assign MEM[48463] = MEM[47060] + MEM[47112];
assign MEM[48464] = MEM[47061] + MEM[47141];
assign MEM[48465] = MEM[47062] + MEM[47136];
assign MEM[48466] = MEM[47063] + MEM[47133];
assign MEM[48467] = MEM[47064] + MEM[47131];
assign MEM[48468] = MEM[47067] + MEM[47171];
assign MEM[48469] = MEM[47069] + MEM[47143];
assign MEM[48470] = MEM[47070] + MEM[47120];
assign MEM[48471] = MEM[47071] + MEM[47138];
assign MEM[48472] = MEM[47074] + MEM[47134];
assign MEM[48473] = MEM[47075] + MEM[47173];
assign MEM[48474] = MEM[47077] + MEM[47150];
assign MEM[48475] = MEM[47080] + MEM[47160];
assign MEM[48476] = MEM[47084] + MEM[47117];
assign MEM[48477] = MEM[47085] + MEM[47154];
assign MEM[48478] = MEM[47087] + MEM[47153];
assign MEM[48479] = MEM[47089] + MEM[47135];
assign MEM[48480] = MEM[47091] + MEM[47139];
assign MEM[48481] = MEM[47093] + MEM[47146];
assign MEM[48482] = MEM[47094] + MEM[47149];
assign MEM[48483] = MEM[47095] + MEM[47205];
assign MEM[48484] = MEM[47096] + MEM[47137];
assign MEM[48485] = MEM[47097] + MEM[47220];
assign MEM[48486] = MEM[47098] + MEM[47157];
assign MEM[48487] = MEM[47099] + MEM[47132];
assign MEM[48488] = MEM[47101] + MEM[47142];
assign MEM[48489] = MEM[47103] + MEM[47147];
assign MEM[48490] = MEM[47104] + MEM[47172];
assign MEM[48491] = MEM[47105] + MEM[47201];
assign MEM[48492] = MEM[47110] + MEM[47185];
assign MEM[48493] = MEM[47113] + MEM[47189];
assign MEM[48494] = MEM[47116] + MEM[47161];
assign MEM[48495] = MEM[47118] + MEM[47208];
assign MEM[48496] = MEM[47119] + MEM[47166];
assign MEM[48497] = MEM[47122] + MEM[47158];
assign MEM[48498] = MEM[47123] + MEM[47183];
assign MEM[48499] = MEM[47124] + MEM[47182];
assign MEM[48500] = MEM[47128] + MEM[47177];
assign MEM[48501] = MEM[47130] + MEM[47186];
assign MEM[48502] = MEM[47140] + MEM[47181];
assign MEM[48503] = MEM[47145] + MEM[47197];
assign MEM[48504] = MEM[47151] + MEM[47241];
assign MEM[48505] = MEM[47152] + MEM[47211];
assign MEM[48506] = MEM[47155] + MEM[47209];
assign MEM[48507] = MEM[47156] + MEM[47195];
assign MEM[48508] = MEM[47159] + MEM[47263];
assign MEM[48509] = MEM[47162] + MEM[47236];
assign MEM[48510] = MEM[47163] + MEM[47230];
assign MEM[48511] = MEM[47164] + MEM[47228];
assign MEM[48512] = MEM[47165] + MEM[47226];
assign MEM[48513] = MEM[47167] + MEM[47229];
assign MEM[48514] = MEM[47168] + MEM[47210];
assign MEM[48515] = MEM[47169] + MEM[47242];
assign MEM[48516] = MEM[47170] + MEM[47221];
assign MEM[48517] = MEM[47174] + MEM[47249];
assign MEM[48518] = MEM[47175] + MEM[47243];
assign MEM[48519] = MEM[47176] + MEM[47267];
assign MEM[48520] = MEM[47178] + MEM[47222];
assign MEM[48521] = MEM[47179] + MEM[47227];
assign MEM[48522] = MEM[47180] + MEM[47256];
assign MEM[48523] = MEM[47184] + MEM[47240];
assign MEM[48524] = MEM[47187] + MEM[47265];
assign MEM[48525] = MEM[47188] + MEM[47266];
assign MEM[48526] = MEM[47190] + MEM[47269];
assign MEM[48527] = MEM[47191] + MEM[47231];
assign MEM[48528] = MEM[47192] + MEM[47289];
assign MEM[48529] = MEM[47193] + MEM[47262];
assign MEM[48530] = MEM[47194] + MEM[47272];
assign MEM[48531] = MEM[47196] + MEM[47253];
assign MEM[48532] = MEM[47198] + MEM[47276];
assign MEM[48533] = MEM[47199] + MEM[47251];
assign MEM[48534] = MEM[47200] + MEM[47270];
assign MEM[48535] = MEM[47202] + MEM[47255];
assign MEM[48536] = MEM[47203] + MEM[47274];
assign MEM[48537] = MEM[47204] + MEM[47257];
assign MEM[48538] = MEM[47206] + MEM[47237];
assign MEM[48539] = MEM[47207] + MEM[47346];
assign MEM[48540] = MEM[47212] + MEM[47309];
assign MEM[48541] = MEM[47213] + MEM[47280];
assign MEM[48542] = MEM[47214] + MEM[47288];
assign MEM[48543] = MEM[47215] + MEM[47295];
assign MEM[48544] = MEM[47216] + MEM[47245];
assign MEM[48545] = MEM[47217] + MEM[47278];
assign MEM[48546] = MEM[47218] + MEM[47300];
assign MEM[48547] = MEM[47219] + MEM[47287];
assign MEM[48548] = MEM[47223] + MEM[47277];
assign MEM[48549] = MEM[47224] + MEM[47291];
assign MEM[48550] = MEM[47225] + MEM[47307];
assign MEM[48551] = MEM[47232] + MEM[47294];
assign MEM[48552] = MEM[47233] + MEM[47279];
assign MEM[48553] = MEM[47234] + MEM[47281];
assign MEM[48554] = MEM[47235] + MEM[47273];
assign MEM[48555] = MEM[47238] + MEM[47301];
assign MEM[48556] = MEM[47239] + MEM[47292];
assign MEM[48557] = MEM[47244] + MEM[47311];
assign MEM[48558] = MEM[47246] + MEM[47302];
assign MEM[48559] = MEM[47247] + MEM[47303];
assign MEM[48560] = MEM[47248] + MEM[47296];
assign MEM[48561] = MEM[47250] + MEM[47316];
assign MEM[48562] = MEM[47252] + MEM[47351];
assign MEM[48563] = MEM[47254] + MEM[47310];
assign MEM[48564] = MEM[47258] + MEM[47336];
assign MEM[48565] = MEM[47259] + MEM[47329];
assign MEM[48566] = MEM[47260] + MEM[47360];
assign MEM[48567] = MEM[47261] + MEM[47335];
assign MEM[48568] = MEM[47264] + MEM[47342];
assign MEM[48569] = MEM[47268] + MEM[47332];
assign MEM[48570] = MEM[47271] + MEM[47352];
assign MEM[48571] = MEM[47275] + MEM[47330];
assign MEM[48572] = MEM[47282] + MEM[47347];
assign MEM[48573] = MEM[47283] + MEM[47322];
assign MEM[48574] = MEM[47284] + MEM[47385];
assign MEM[48575] = MEM[47285] + MEM[47355];
assign MEM[48576] = MEM[47286] + MEM[47317];
assign MEM[48577] = MEM[47290] + MEM[47345];
assign MEM[48578] = MEM[47293] + MEM[47410];
assign MEM[48579] = MEM[47297] + MEM[47371];
assign MEM[48580] = MEM[47298] + MEM[47359];
assign MEM[48581] = MEM[47299] + MEM[47354];
assign MEM[48582] = MEM[47304] + MEM[47340];
assign MEM[48583] = MEM[47305] + MEM[47356];
assign MEM[48584] = MEM[47306] + MEM[47337];
assign MEM[48585] = MEM[47308] + MEM[47390];
assign MEM[48586] = MEM[47312] + MEM[47396];
assign MEM[48587] = MEM[47313] + MEM[47367];
assign MEM[48588] = MEM[47314] + MEM[47393];
assign MEM[48589] = MEM[47315] + MEM[47387];
assign MEM[48590] = MEM[47318] + MEM[47397];
assign MEM[48591] = MEM[47319] + MEM[47363];
assign MEM[48592] = MEM[47320] + MEM[47399];
assign MEM[48593] = MEM[47321] + MEM[47349];
assign MEM[48594] = MEM[47323] + MEM[47413];
assign MEM[48595] = MEM[47324] + MEM[47372];
assign MEM[48596] = MEM[47325] + MEM[47408];
assign MEM[48597] = MEM[47326] + MEM[47428];
assign MEM[48598] = MEM[47327] + MEM[47378];
assign MEM[48599] = MEM[47328] + MEM[47405];
assign MEM[48600] = MEM[47331] + MEM[47374];
assign MEM[48601] = MEM[47333] + MEM[47392];
assign MEM[48602] = MEM[47334] + MEM[47394];
assign MEM[48603] = MEM[47338] + MEM[47409];
assign MEM[48604] = MEM[47339] + MEM[47380];
assign MEM[48605] = MEM[47341] + MEM[47384];
assign MEM[48606] = MEM[47343] + MEM[47401];
assign MEM[48607] = MEM[47344] + MEM[47388];
assign MEM[48608] = MEM[47348] + MEM[47418];
assign MEM[48609] = MEM[47350] + MEM[47400];
assign MEM[48610] = MEM[47353] + MEM[47419];
assign MEM[48611] = MEM[47357] + MEM[47411];
assign MEM[48612] = MEM[47358] + MEM[47398];
assign MEM[48613] = MEM[47361] + MEM[47412];
assign MEM[48614] = MEM[47362] + MEM[47488];
assign MEM[48615] = MEM[47364] + MEM[47433];
assign MEM[48616] = MEM[47365] + MEM[47417];
assign MEM[48617] = MEM[47366] + MEM[47420];
assign MEM[48618] = MEM[47368] + MEM[47415];
assign MEM[48619] = MEM[47369] + MEM[47426];
assign MEM[48620] = MEM[47370] + MEM[47440];
assign MEM[48621] = MEM[47373] + MEM[47447];
assign MEM[48622] = MEM[47375] + MEM[47439];
assign MEM[48623] = MEM[47376] + MEM[47423];
assign MEM[48624] = MEM[47377] + MEM[47431];
assign MEM[48625] = MEM[47379] + MEM[47462];
assign MEM[48626] = MEM[47381] + MEM[47429];
assign MEM[48627] = MEM[47382] + MEM[47450];
assign MEM[48628] = MEM[47383] + MEM[47465];
assign MEM[48629] = MEM[47386] + MEM[47461];
assign MEM[48630] = MEM[47389] + MEM[47432];
assign MEM[48631] = MEM[47391] + MEM[47464];
assign MEM[48632] = MEM[47395] + MEM[47476];
assign MEM[48633] = MEM[47402] + MEM[47457];
assign MEM[48634] = MEM[47403] + MEM[47444];
assign MEM[48635] = MEM[47404] + MEM[47487];
assign MEM[48636] = MEM[47406] + MEM[47454];
assign MEM[48637] = MEM[47407] + MEM[47458];
assign MEM[48638] = MEM[47414] + MEM[47483];
assign MEM[48639] = MEM[47416] + MEM[47451];
assign MEM[48640] = MEM[47421] + MEM[47491];
assign MEM[48641] = MEM[47422] + MEM[47470];
assign MEM[48642] = MEM[47424] + MEM[47489];
assign MEM[48643] = MEM[47425] + MEM[47547];
assign MEM[48644] = MEM[47427] + MEM[47482];
assign MEM[48645] = MEM[47430] + MEM[47478];
assign MEM[48646] = MEM[47434] + MEM[47493];
assign MEM[48647] = MEM[47435] + MEM[47512];
assign MEM[48648] = MEM[47436] + MEM[47504];
assign MEM[48649] = MEM[47437] + MEM[47513];
assign MEM[48650] = MEM[47438] + MEM[47497];
assign MEM[48651] = MEM[47441] + MEM[47485];
assign MEM[48652] = MEM[47442] + MEM[47498];
assign MEM[48653] = MEM[47443] + MEM[47506];
assign MEM[48654] = MEM[47445] + MEM[47518];
assign MEM[48655] = MEM[47446] + MEM[47519];
assign MEM[48656] = MEM[47448] + MEM[47516];
assign MEM[48657] = MEM[47449] + MEM[47511];
assign MEM[48658] = MEM[47452] + MEM[47530];
assign MEM[48659] = MEM[47453] + MEM[47532];
assign MEM[48660] = MEM[47455] + MEM[47514];
assign MEM[48661] = MEM[47456] + MEM[47515];
assign MEM[48662] = MEM[47459] + MEM[47520];
assign MEM[48663] = MEM[47460] + MEM[47559];
assign MEM[48664] = MEM[47463] + MEM[47505];
assign MEM[48665] = MEM[47466] + MEM[47529];
assign MEM[48666] = MEM[47467] + MEM[47556];
assign MEM[48667] = MEM[47468] + MEM[47521];
assign MEM[48668] = MEM[47469] + MEM[47536];
assign MEM[48669] = MEM[47471] + MEM[47606];
assign MEM[48670] = MEM[47472] + MEM[47552];
assign MEM[48671] = MEM[47473] + MEM[47535];
assign MEM[48672] = MEM[47474] + MEM[47548];
assign MEM[48673] = MEM[47475] + MEM[47551];
assign MEM[48674] = MEM[47477] + MEM[47558];
assign MEM[48675] = MEM[47479] + MEM[47524];
assign MEM[48676] = MEM[47480] + MEM[47537];
assign MEM[48677] = MEM[47481] + MEM[47578];
assign MEM[48678] = MEM[47484] + MEM[47553];
assign MEM[48679] = MEM[47486] + MEM[47526];
assign MEM[48680] = MEM[47490] + MEM[47582];
assign MEM[48681] = MEM[47492] + MEM[47531];
assign MEM[48682] = MEM[47494] + MEM[47545];
assign MEM[48683] = MEM[47495] + MEM[47561];
assign MEM[48684] = MEM[47496] + MEM[47580];
assign MEM[48685] = MEM[47499] + MEM[47549];
assign MEM[48686] = MEM[47500] + MEM[47563];
assign MEM[48687] = MEM[47501] + MEM[47587];
assign MEM[48688] = MEM[47502] + MEM[47554];
assign MEM[48689] = MEM[47503] + MEM[47568];
assign MEM[48690] = MEM[47507] + MEM[47575];
assign MEM[48691] = MEM[47508] + MEM[47614];
assign MEM[48692] = MEM[47509] + MEM[47539];
assign MEM[48693] = MEM[47510] + MEM[47571];
assign MEM[48694] = MEM[47517] + MEM[47565];
assign MEM[48695] = MEM[47522] + MEM[47555];
assign MEM[48696] = MEM[47523] + MEM[47570];
assign MEM[48697] = MEM[47525] + MEM[47610];
assign MEM[48698] = MEM[47527] + MEM[47609];
assign MEM[48699] = MEM[47528] + MEM[47618];
assign MEM[48700] = MEM[47533] + MEM[47589];
assign MEM[48701] = MEM[47534] + MEM[47605];
assign MEM[48702] = MEM[47538] + MEM[47648];
assign MEM[48703] = MEM[47540] + MEM[47569];
assign MEM[48704] = MEM[47541] + MEM[47647];
assign MEM[48705] = MEM[47542] + MEM[47600];
assign MEM[48706] = MEM[47543] + MEM[47622];
assign MEM[48707] = MEM[47544] + MEM[47595];
assign MEM[48708] = MEM[47546] + MEM[47584];
assign MEM[48709] = MEM[47550] + MEM[47583];
assign MEM[48710] = MEM[47557] + MEM[47615];
assign MEM[48711] = MEM[47560] + MEM[47626];
assign MEM[48712] = MEM[47562] + MEM[47656];
assign MEM[48713] = MEM[47564] + MEM[47627];
assign MEM[48714] = MEM[47566] + MEM[47658];
assign MEM[48715] = MEM[47567] + MEM[47599];
assign MEM[48716] = MEM[47572] + MEM[47651];
assign MEM[48717] = MEM[47573] + MEM[47633];
assign MEM[48718] = MEM[47574] + MEM[47636];
assign MEM[48719] = MEM[47576] + MEM[47687];
assign MEM[48720] = MEM[47577] + MEM[47628];
assign MEM[48721] = MEM[47579] + MEM[47632];
assign MEM[48722] = MEM[47581] + MEM[47643];
assign MEM[48723] = MEM[47585] + MEM[47638];
assign MEM[48724] = MEM[47586] + MEM[47661];
assign MEM[48725] = MEM[47588] + MEM[47660];
assign MEM[48726] = MEM[47590] + MEM[47677];
assign MEM[48727] = MEM[47591] + MEM[47649];
assign MEM[48728] = MEM[47592] + MEM[47640];
assign MEM[48729] = MEM[47593] + MEM[47637];
assign MEM[48730] = MEM[47594] + MEM[47672];
assign MEM[48731] = MEM[47596] + MEM[47652];
assign MEM[48732] = MEM[47597] + MEM[47653];
assign MEM[48733] = MEM[47598] + MEM[47666];
assign MEM[48734] = MEM[47601] + MEM[47673];
assign MEM[48735] = MEM[47602] + MEM[47662];
assign MEM[48736] = MEM[47603] + MEM[47680];
assign MEM[48737] = MEM[47604] + MEM[47645];
assign MEM[48738] = MEM[47607] + MEM[47671];
assign MEM[48739] = MEM[47608] + MEM[47668];
assign MEM[48740] = MEM[47611] + MEM[47644];
assign MEM[48741] = MEM[47612] + MEM[47681];
assign MEM[48742] = MEM[47613] + MEM[47657];
assign MEM[48743] = MEM[47616] + MEM[47678];
assign MEM[48744] = MEM[47617] + MEM[47634];
assign MEM[48745] = MEM[47619] + MEM[47695];
assign MEM[48746] = MEM[47620] + MEM[47691];
assign MEM[48747] = MEM[47621] + MEM[47699];
assign MEM[48748] = MEM[47623] + MEM[47697];
assign MEM[48749] = MEM[47624] + MEM[47692];
assign MEM[48750] = MEM[47625] + MEM[47683];
assign MEM[48751] = MEM[47629] + MEM[47667];
assign MEM[48752] = MEM[47630] + MEM[47686];
assign MEM[48753] = MEM[47631] + MEM[47756];
assign MEM[48754] = MEM[47635] + MEM[47694];
assign MEM[48755] = MEM[47639] + MEM[47679];
assign MEM[48756] = MEM[47641] + MEM[47722];
assign MEM[48757] = MEM[47642] + MEM[47701];
assign MEM[48758] = MEM[47646] + MEM[47709];
assign MEM[48759] = MEM[47650] + MEM[47698];
assign MEM[48760] = MEM[47654] + MEM[47718];
assign MEM[48761] = MEM[47655] + MEM[47704];
assign MEM[48762] = MEM[47659] + MEM[47711];
assign MEM[48763] = MEM[47663] + MEM[47746];
assign MEM[48764] = MEM[47664] + MEM[47714];
assign MEM[48765] = MEM[47665] + MEM[47736];
assign MEM[48766] = MEM[47669] + MEM[47745];
assign MEM[48767] = MEM[47670] + MEM[47787];
assign MEM[48768] = MEM[47674] + MEM[47729];
assign MEM[48769] = MEM[47675] + MEM[47752];
assign MEM[48770] = MEM[47676] + MEM[47728];
assign MEM[48771] = MEM[47682] + MEM[47735];
assign MEM[48772] = MEM[47684] + MEM[47772];
assign MEM[48773] = MEM[47685] + MEM[47739];
assign MEM[48774] = MEM[47688] + MEM[47761];
assign MEM[48775] = MEM[47689] + MEM[47785];
assign MEM[48776] = MEM[47690] + MEM[47751];
assign MEM[48777] = MEM[47693] + MEM[47760];
assign MEM[48778] = MEM[47696] + MEM[47776];
assign MEM[48779] = MEM[47700] + MEM[47754];
assign MEM[48780] = MEM[47702] + MEM[47784];
assign MEM[48781] = MEM[47703] + MEM[47793];
assign MEM[48782] = MEM[47705] + MEM[47768];
assign MEM[48783] = MEM[47706] + MEM[47782];
assign MEM[48784] = MEM[47707] + MEM[47764];
assign MEM[48785] = MEM[47708] + MEM[47741];
assign MEM[48786] = MEM[47710] + MEM[47771];
assign MEM[48787] = MEM[47712] + MEM[47794];
assign MEM[48788] = MEM[47713] + MEM[47781];
assign MEM[48789] = MEM[47715] + MEM[47791];
assign MEM[48790] = MEM[47716] + MEM[47744];
assign MEM[48791] = MEM[47717] + MEM[47778];
assign MEM[48792] = MEM[47719] + MEM[47815];
assign MEM[48793] = MEM[47720] + MEM[47786];
assign MEM[48794] = MEM[47721] + MEM[47773];
assign MEM[48795] = MEM[47723] + MEM[47779];
assign MEM[48796] = MEM[47724] + MEM[47769];
assign MEM[48797] = MEM[47725] + MEM[47770];
assign MEM[48798] = MEM[47726] + MEM[47795];
assign MEM[48799] = MEM[47727] + MEM[47758];
assign MEM[48800] = MEM[47730] + MEM[47797];
assign MEM[48801] = MEM[47731] + MEM[47800];
assign MEM[48802] = MEM[47732] + MEM[47775];
assign MEM[48803] = MEM[47733] + MEM[47790];
assign MEM[48804] = MEM[47734] + MEM[47767];
assign MEM[48805] = MEM[47737] + MEM[47806];
assign MEM[48806] = MEM[47738] + MEM[47805];
assign MEM[48807] = MEM[47740] + MEM[47789];
assign MEM[48808] = MEM[47742] + MEM[47812];
assign MEM[48809] = MEM[47743] + MEM[47829];
assign MEM[48810] = MEM[47747] + MEM[47809];
assign MEM[48811] = MEM[47748] + MEM[47860];
assign MEM[48812] = MEM[47749] + MEM[47838];
assign MEM[48813] = MEM[47750] + MEM[47844];
assign MEM[48814] = MEM[47753] + MEM[47826];
assign MEM[48815] = MEM[47755] + MEM[47832];
assign MEM[48816] = MEM[47757] + MEM[47801];
assign MEM[48817] = MEM[47759] + MEM[47822];
assign MEM[48818] = MEM[47762] + MEM[47867];
assign MEM[48819] = MEM[47763] + MEM[47803];
assign MEM[48820] = MEM[47765] + MEM[47847];
assign MEM[48821] = MEM[47766] + MEM[47825];
assign MEM[48822] = MEM[47774] + MEM[47802];
assign MEM[48823] = MEM[47777] + MEM[47841];
assign MEM[48824] = MEM[47780] + MEM[47818];
assign MEM[48825] = MEM[47783] + MEM[47819];
assign MEM[48826] = MEM[47788] + MEM[47853];
assign MEM[48827] = MEM[47792] + MEM[47870];
assign MEM[48828] = MEM[47796] + MEM[47859];
assign MEM[48829] = MEM[47798] + MEM[47878];
assign MEM[48830] = MEM[47799] + MEM[47854];
assign MEM[48831] = MEM[47804] + MEM[47888];
assign MEM[48832] = MEM[47807] + MEM[47851];
assign MEM[48833] = MEM[47808] + MEM[47876];
assign MEM[48834] = MEM[47810] + MEM[47917];
assign MEM[48835] = MEM[47811] + MEM[47856];
assign MEM[48836] = MEM[47813] + MEM[47873];
assign MEM[48837] = MEM[47814] + MEM[47874];
assign MEM[48838] = MEM[47816] + MEM[47849];
assign MEM[48839] = MEM[47817] + MEM[47882];
assign MEM[48840] = MEM[47820] + MEM[47905];
assign MEM[48841] = MEM[47821] + MEM[47891];
assign MEM[48842] = MEM[47823] + MEM[47896];
assign MEM[48843] = MEM[47824] + MEM[47913];
assign MEM[48844] = MEM[47827] + MEM[47919];
assign MEM[48845] = MEM[47828] + MEM[47898];
assign MEM[48846] = MEM[47830] + MEM[47900];
assign MEM[48847] = MEM[47831] + MEM[47921];
assign MEM[48848] = MEM[47833] + MEM[47911];
assign MEM[48849] = MEM[47834] + MEM[47865];
assign MEM[48850] = MEM[47835] + MEM[47909];
assign MEM[48851] = MEM[47836] + MEM[47877];
assign MEM[48852] = MEM[47837] + MEM[47883];
assign MEM[48853] = MEM[47839] + MEM[47886];
assign MEM[48854] = MEM[47840] + MEM[47920];
assign MEM[48855] = MEM[47842] + MEM[47906];
assign MEM[48856] = MEM[47843] + MEM[47910];
assign MEM[48857] = MEM[47845] + MEM[47902];
assign MEM[48858] = MEM[47846] + MEM[47864];
assign MEM[48859] = MEM[47848] + MEM[47887];
assign MEM[48860] = MEM[47850] + MEM[47912];
assign MEM[48861] = MEM[47852] + MEM[47914];
assign MEM[48862] = MEM[47855] + MEM[47922];
assign MEM[48863] = MEM[47857] + MEM[47885];
assign MEM[48864] = MEM[47858] + MEM[47916];
assign MEM[48865] = MEM[47861] + MEM[47908];
assign MEM[48866] = MEM[47862] + MEM[47934];
assign MEM[48867] = MEM[47863] + MEM[47960];
assign MEM[48868] = MEM[47866] + MEM[47954];
assign MEM[48869] = MEM[47868] + MEM[47945];
assign MEM[48870] = MEM[47869] + MEM[47928];
assign MEM[48871] = MEM[47871] + MEM[47938];
assign MEM[48872] = MEM[47872] + MEM[47927];
assign MEM[48873] = MEM[47875] + MEM[47959];
assign MEM[48874] = MEM[47879] + MEM[47918];
assign MEM[48875] = MEM[47880] + MEM[47925];
assign MEM[48876] = MEM[47881] + MEM[47931];
assign MEM[48877] = MEM[47884] + MEM[47965];
assign MEM[48878] = MEM[47889] + MEM[47987];
assign MEM[48879] = MEM[47890] + MEM[47941];
assign MEM[48880] = MEM[47892] + MEM[47967];
assign MEM[48881] = MEM[47893] + MEM[47984];
assign MEM[48882] = MEM[47894] + MEM[47991];
assign MEM[48883] = MEM[47895] + MEM[47944];
assign MEM[48884] = MEM[47897] + MEM[47948];
assign MEM[48885] = MEM[47899] + MEM[47988];
assign MEM[48886] = MEM[47901] + MEM[47973];
assign MEM[48887] = MEM[47903] + MEM[47969];
assign MEM[48888] = MEM[47904] + MEM[47958];
assign MEM[48889] = MEM[47907] + MEM[47995];
assign MEM[48890] = MEM[47915] + MEM[47979];
assign MEM[48891] = MEM[47923] + MEM[47974];
assign MEM[48892] = MEM[47924] + MEM[47975];
assign MEM[48893] = MEM[47926] + MEM[47968];
assign MEM[48894] = MEM[47929] + MEM[47977];
assign MEM[48895] = MEM[47930] + MEM[48016];
assign MEM[48896] = MEM[47932] + MEM[48004];
assign MEM[48897] = MEM[47933] + MEM[47985];
assign MEM[48898] = MEM[47935] + MEM[48010];
assign MEM[48899] = MEM[47936] + MEM[48057];
assign MEM[48900] = MEM[47937] + MEM[47993];
assign MEM[48901] = MEM[47939] + MEM[48025];
assign MEM[48902] = MEM[47940] + MEM[48006];
assign MEM[48903] = MEM[47942] + MEM[48012];
assign MEM[48904] = MEM[47943] + MEM[48007];
assign MEM[48905] = MEM[47946] + MEM[48002];
assign MEM[48906] = MEM[47947] + MEM[47998];
assign MEM[48907] = MEM[47949] + MEM[48011];
assign MEM[48908] = MEM[47950] + MEM[48001];
assign MEM[48909] = MEM[47951] + MEM[48014];
assign MEM[48910] = MEM[47952] + MEM[48000];
assign MEM[48911] = MEM[47953] + MEM[47983];
assign MEM[48912] = MEM[47955] + MEM[48022];
assign MEM[48913] = MEM[47956] + MEM[48031];
assign MEM[48914] = MEM[47957] + MEM[47999];
assign MEM[48915] = MEM[47961] + MEM[48038];
assign MEM[48916] = MEM[47962] + MEM[48061];
assign MEM[48917] = MEM[47963] + MEM[48024];
assign MEM[48918] = MEM[47964] + MEM[48021];
assign MEM[48919] = MEM[47966] + MEM[48029];
assign MEM[48920] = MEM[47970] + MEM[48032];
assign MEM[48921] = MEM[47971] + MEM[48026];
assign MEM[48922] = MEM[47972] + MEM[48070];
assign MEM[48923] = MEM[47976] + MEM[48027];
assign MEM[48924] = MEM[47978] + MEM[48068];
assign MEM[48925] = MEM[47980] + MEM[48023];
assign MEM[48926] = MEM[47981] + MEM[48042];
assign MEM[48927] = MEM[47982] + MEM[48034];
assign MEM[48928] = MEM[47986] + MEM[48043];
assign MEM[48929] = MEM[47989] + MEM[48049];
assign MEM[48930] = MEM[47990] + MEM[48066];
assign MEM[48931] = MEM[47992] + MEM[48064];
assign MEM[48932] = MEM[47994] + MEM[48069];
assign MEM[48933] = MEM[47996] + MEM[48084];
assign MEM[48934] = MEM[47997] + MEM[48055];
assign MEM[48935] = MEM[48003] + MEM[48056];
assign MEM[48936] = MEM[48005] + MEM[48081];
assign MEM[48937] = MEM[48008] + MEM[48104];
assign MEM[48938] = MEM[48009] + MEM[48080];
assign MEM[48939] = MEM[48013] + MEM[48075];
assign MEM[48940] = MEM[48015] + MEM[48077];
assign MEM[48941] = MEM[48017] + MEM[48122];
assign MEM[48942] = MEM[48018] + MEM[48074];
assign MEM[48943] = MEM[48019] + MEM[48082];
assign MEM[48944] = MEM[48020] + MEM[48076];
assign MEM[48945] = MEM[48028] + MEM[48095];
assign MEM[48946] = MEM[48030] + MEM[48101];
assign MEM[48947] = MEM[48033] + MEM[48096];
assign MEM[48948] = MEM[48035] + MEM[48093];
assign MEM[48949] = MEM[48036] + MEM[48098];
assign MEM[48950] = MEM[48037] + MEM[48103];
assign MEM[48951] = MEM[48039] + MEM[48091];
assign MEM[48952] = MEM[48040] + MEM[48107];
assign MEM[48953] = MEM[48041] + MEM[48097];
assign MEM[48954] = MEM[48044] + MEM[48111];
assign MEM[48955] = MEM[48045] + MEM[48105];
assign MEM[48956] = MEM[48046] + MEM[48079];
assign MEM[48957] = MEM[48047] + MEM[48135];
assign MEM[48958] = MEM[48048] + MEM[48133];
assign MEM[48959] = MEM[48050] + MEM[48108];
assign MEM[48960] = MEM[48051] + MEM[48114];
assign MEM[48961] = MEM[48052] + MEM[48106];
assign MEM[48962] = MEM[48053] + MEM[48138];
assign MEM[48963] = MEM[48054] + MEM[48102];
assign MEM[48964] = MEM[48058] + MEM[48162];
assign MEM[48965] = MEM[48059] + MEM[48112];
assign MEM[48966] = MEM[48060] + MEM[48141];
assign MEM[48967] = MEM[48062] + MEM[48115];
assign MEM[48968] = MEM[48063] + MEM[48131];
assign MEM[48969] = MEM[48065] + MEM[48143];
assign MEM[48970] = MEM[48067] + MEM[48121];
assign MEM[48971] = MEM[48071] + MEM[48120];
assign MEM[48972] = MEM[48072] + MEM[48157];
assign MEM[48973] = MEM[48073] + MEM[48150];
assign MEM[48974] = MEM[48078] + MEM[48145];
assign MEM[48975] = MEM[48083] + MEM[48129];
assign MEM[48976] = MEM[48085] + MEM[48165];
assign MEM[48977] = MEM[48086] + MEM[48130];
assign MEM[48978] = MEM[48087] + MEM[48136];
assign MEM[48979] = MEM[48088] + MEM[48147];
assign MEM[48980] = MEM[48089] + MEM[48153];
assign MEM[48981] = MEM[48090] + MEM[48137];
assign MEM[48982] = MEM[48092] + MEM[48142];
assign MEM[48983] = MEM[48094] + MEM[48140];
assign MEM[48984] = MEM[48099] + MEM[48159];
assign MEM[48985] = MEM[48100] + MEM[48148];
assign MEM[48986] = MEM[48109] + MEM[48167];
assign MEM[48987] = MEM[48110] + MEM[48173];
assign MEM[48988] = MEM[48113] + MEM[48193];
assign MEM[48989] = MEM[48116] + MEM[48168];
assign MEM[48990] = MEM[48117] + MEM[48206];
assign MEM[48991] = MEM[48118] + MEM[48211];
assign MEM[48992] = MEM[48119] + MEM[48172];
assign MEM[48993] = MEM[48123] + MEM[48184];
assign MEM[48994] = MEM[48124] + MEM[48198];
assign MEM[48995] = MEM[48125] + MEM[48203];
assign MEM[48996] = MEM[48126] + MEM[48192];
assign MEM[48997] = MEM[48127] + MEM[48181];
assign MEM[48998] = MEM[48128] + MEM[48197];
assign MEM[48999] = MEM[48132] + MEM[48191];
assign MEM[49000] = MEM[48134] + MEM[48209];
assign MEM[49001] = MEM[48139] + MEM[48187];
assign MEM[49002] = MEM[48144] + MEM[48220];
assign MEM[49003] = MEM[48146] + MEM[48183];
assign MEM[49004] = MEM[48149] + MEM[48213];
assign MEM[49005] = MEM[48151] + MEM[48217];
assign MEM[49006] = MEM[48152] + MEM[48223];
assign MEM[49007] = MEM[48154] + MEM[48228];
assign MEM[49008] = MEM[48155] + MEM[48218];
assign MEM[49009] = MEM[48156] + MEM[48196];
assign MEM[49010] = MEM[48158] + MEM[48248];
assign MEM[49011] = MEM[48160] + MEM[48210];
assign MEM[49012] = MEM[48161] + MEM[48219];
assign MEM[49013] = MEM[48163] + MEM[48239];
assign MEM[49014] = MEM[48164] + MEM[48255];
assign MEM[49015] = MEM[48166] + MEM[48205];
assign MEM[49016] = MEM[48169] + MEM[48236];
assign MEM[49017] = MEM[48170] + MEM[48216];
assign MEM[49018] = MEM[48171] + MEM[48247];
assign MEM[49019] = MEM[48174] + MEM[48226];
assign MEM[49020] = MEM[48175] + MEM[48257];
assign MEM[49021] = MEM[48176] + MEM[48232];
assign MEM[49022] = MEM[48177] + MEM[48234];
assign MEM[49023] = MEM[48178] + MEM[48258];
assign MEM[49024] = MEM[48179] + MEM[48272];
assign MEM[49025] = MEM[48180] + MEM[48238];
assign MEM[49026] = MEM[48182] + MEM[48222];
assign MEM[49027] = MEM[48185] + MEM[48229];
assign MEM[49028] = MEM[48186] + MEM[48235];
assign MEM[49029] = MEM[48188] + MEM[48265];
assign MEM[49030] = MEM[48189] + MEM[48260];
assign MEM[49031] = MEM[48190] + MEM[48280];
assign MEM[49032] = MEM[48194] + MEM[48268];
assign MEM[49033] = MEM[48195] + MEM[48253];
assign MEM[49034] = MEM[48199] + MEM[48249];
assign MEM[49035] = MEM[48200] + MEM[48246];
assign MEM[49036] = MEM[48201] + MEM[48250];
assign MEM[49037] = MEM[48202] + MEM[48244];
assign MEM[49038] = MEM[48204] + MEM[48245];
assign MEM[49039] = MEM[48207] + MEM[48251];
assign MEM[49040] = MEM[48208] + MEM[48281];
assign MEM[49041] = MEM[48212] + MEM[48285];
assign MEM[49042] = MEM[48214] + MEM[48274];
assign MEM[49043] = MEM[48215] + MEM[48313];
assign MEM[49044] = MEM[48221] + MEM[48294];
assign MEM[49045] = MEM[48224] + MEM[48302];
assign MEM[49046] = MEM[48225] + MEM[48291];
assign MEM[49047] = MEM[48227] + MEM[48286];
assign MEM[49048] = MEM[48230] + MEM[48310];
assign MEM[49049] = MEM[48231] + MEM[48306];
assign MEM[49050] = MEM[48233] + MEM[48304];
assign MEM[49051] = MEM[48237] + MEM[48292];
assign MEM[49052] = MEM[48240] + MEM[48324];
assign MEM[49053] = MEM[48241] + MEM[48326];
assign MEM[49054] = MEM[48242] + MEM[48314];
assign MEM[49055] = MEM[48243] + MEM[48329];
assign MEM[49056] = MEM[48252] + MEM[48301];
assign MEM[49057] = MEM[48254] + MEM[48312];
assign MEM[49058] = MEM[48256] + MEM[48299];
assign MEM[49059] = MEM[48259] + MEM[48357];
assign MEM[49060] = MEM[48261] + MEM[48330];
assign MEM[49061] = MEM[48262] + MEM[48323];
assign MEM[49062] = MEM[48263] + MEM[48315];
assign MEM[49063] = MEM[48264] + MEM[48322];
assign MEM[49064] = MEM[48266] + MEM[48289];
assign MEM[49065] = MEM[48267] + MEM[48316];
assign MEM[49066] = MEM[48269] + MEM[48334];
assign MEM[49067] = MEM[48270] + MEM[48335];
assign MEM[49068] = MEM[48271] + MEM[48340];
assign MEM[49069] = MEM[48273] + MEM[48297];
assign MEM[49070] = MEM[48275] + MEM[48331];
assign MEM[49071] = MEM[48276] + MEM[48341];
assign MEM[49072] = MEM[48277] + MEM[48351];
assign MEM[49073] = MEM[48278] + MEM[48394];
assign MEM[49074] = MEM[48279] + MEM[48373];
assign MEM[49075] = MEM[48282] + MEM[48336];
assign MEM[49076] = MEM[48283] + MEM[48348];
assign MEM[49077] = MEM[48284] + MEM[48395];
assign MEM[49078] = MEM[48287] + MEM[48343];
assign MEM[49079] = MEM[48288] + MEM[48372];
assign MEM[49080] = MEM[48290] + MEM[48356];
assign MEM[49081] = MEM[48293] + MEM[48370];
assign MEM[49082] = MEM[48295] + MEM[48378];
assign MEM[49083] = MEM[48296] + MEM[48342];
assign MEM[49084] = MEM[48298] + MEM[48344];
assign MEM[49085] = MEM[48300] + MEM[48383];
assign MEM[49086] = MEM[48303] + MEM[48362];
assign MEM[49087] = MEM[48305] + MEM[48375];
assign MEM[49088] = MEM[48307] + MEM[48387];
assign MEM[49089] = MEM[48308] + MEM[48365];
assign MEM[49090] = MEM[48309] + MEM[48376];
assign MEM[49091] = MEM[48311] + MEM[48374];
assign MEM[49092] = MEM[48317] + MEM[48367];
assign MEM[49093] = MEM[48318] + MEM[48360];
assign MEM[49094] = MEM[48319] + MEM[48359];
assign MEM[49095] = MEM[48320] + MEM[48381];
assign MEM[49096] = MEM[48321] + MEM[48399];
assign MEM[49097] = MEM[48325] + MEM[48382];
assign MEM[49098] = MEM[48327] + MEM[48400];
assign MEM[49099] = MEM[48328] + MEM[48379];
assign MEM[49100] = MEM[48332] + MEM[48420];
assign MEM[49101] = MEM[48333] + MEM[48401];
assign MEM[49102] = MEM[48337] + MEM[48391];
assign MEM[49103] = MEM[48338] + MEM[48408];
assign MEM[49104] = MEM[48339] + MEM[48386];
assign MEM[49105] = MEM[48345] + MEM[48428];
assign MEM[49106] = MEM[48346] + MEM[48413];
assign MEM[49107] = MEM[48347] + MEM[48416];
assign MEM[49108] = MEM[48349] + MEM[48417];
assign MEM[49109] = MEM[48350] + MEM[48435];
assign MEM[49110] = MEM[48352] + MEM[48409];
assign MEM[49111] = MEM[48353] + MEM[48402];
assign MEM[49112] = MEM[48354] + MEM[48418];
assign MEM[49113] = MEM[48355] + MEM[48412];
assign MEM[49114] = MEM[48358] + MEM[48425];
assign MEM[49115] = MEM[48361] + MEM[48419];
assign MEM[49116] = MEM[48363] + MEM[48426];
assign MEM[49117] = MEM[48364] + MEM[48415];
assign MEM[49118] = MEM[48366] + MEM[48405];
assign MEM[49119] = MEM[48368] + MEM[48441];
assign MEM[49120] = MEM[48369] + MEM[48439];
assign MEM[49121] = MEM[48371] + MEM[48432];
assign MEM[49122] = MEM[48377] + MEM[48472];
assign MEM[49123] = MEM[48380] + MEM[48449];
assign MEM[49124] = MEM[48384] + MEM[48494];
assign MEM[49125] = MEM[48385] + MEM[48453];
assign MEM[49126] = MEM[48388] + MEM[48454];
assign MEM[49127] = MEM[48389] + MEM[48445];
assign MEM[49128] = MEM[48390] + MEM[48440];
assign MEM[49129] = MEM[48392] + MEM[48423];
assign MEM[49130] = MEM[48393] + MEM[48444];
assign MEM[49131] = MEM[48396] + MEM[48473];
assign MEM[49132] = MEM[48397] + MEM[48462];
assign MEM[49133] = MEM[48398] + MEM[48455];
assign MEM[49134] = MEM[48403] + MEM[48471];
assign MEM[49135] = MEM[48404] + MEM[48466];
assign MEM[49136] = MEM[48406] + MEM[48461];
assign MEM[49137] = MEM[48407] + MEM[48470];
assign MEM[49138] = MEM[48410] + MEM[48484];
assign MEM[49139] = MEM[48411] + MEM[48493];
assign MEM[49140] = MEM[48414] + MEM[48476];
assign MEM[49141] = MEM[48421] + MEM[48497];
assign MEM[49142] = MEM[48422] + MEM[48477];
assign MEM[49143] = MEM[48424] + MEM[48500];
assign MEM[49144] = MEM[48427] + MEM[48498];
assign MEM[49145] = MEM[48429] + MEM[48495];
assign MEM[49146] = MEM[48430] + MEM[48483];
assign MEM[49147] = MEM[48431] + MEM[48489];
assign MEM[49148] = MEM[48433] + MEM[48490];
assign MEM[49149] = MEM[48434] + MEM[48474];
assign MEM[49150] = MEM[48436] + MEM[48521];
assign MEM[49151] = MEM[48437] + MEM[48479];
assign MEM[49152] = MEM[48438] + MEM[48504];
assign MEM[49153] = MEM[48442] + MEM[48496];
assign MEM[49154] = MEM[48443] + MEM[48506];
assign MEM[49155] = MEM[48446] + MEM[48532];
assign MEM[49156] = MEM[48447] + MEM[48524];
assign MEM[49157] = MEM[48448] + MEM[48541];
assign MEM[49158] = MEM[48450] + MEM[48499];
assign MEM[49159] = MEM[48451] + MEM[48507];
assign MEM[49160] = MEM[48452] + MEM[48542];
assign MEM[49161] = MEM[48456] + MEM[48534];
assign MEM[49162] = MEM[48457] + MEM[48528];
assign MEM[49163] = MEM[48458] + MEM[48517];
assign MEM[49164] = MEM[48459] + MEM[48508];
assign MEM[49165] = MEM[48460] + MEM[48556];
assign MEM[49166] = MEM[48463] + MEM[48503];
assign MEM[49167] = MEM[48464] + MEM[48525];
assign MEM[49168] = MEM[48465] + MEM[48533];
assign MEM[49169] = MEM[48467] + MEM[48520];
assign MEM[49170] = MEM[48468] + MEM[48557];
assign MEM[49171] = MEM[48469] + MEM[48519];
assign MEM[49172] = MEM[48475] + MEM[48551];
assign MEM[49173] = MEM[48478] + MEM[48578];
assign MEM[49174] = MEM[48480] + MEM[48537];
assign MEM[49175] = MEM[48481] + MEM[48540];
assign MEM[49176] = MEM[48482] + MEM[48543];
assign MEM[49177] = MEM[48485] + MEM[48569];
assign MEM[49178] = MEM[48486] + MEM[48547];
assign MEM[49179] = MEM[48487] + MEM[48535];
assign MEM[49180] = MEM[48488] + MEM[48509];
assign MEM[49181] = MEM[48491] + MEM[48555];
assign MEM[49182] = MEM[48492] + MEM[48560];
assign MEM[49183] = MEM[48501] + MEM[48546];
assign MEM[49184] = MEM[48502] + MEM[48575];
assign MEM[49185] = MEM[48505] + MEM[48564];
assign MEM[49186] = MEM[48510] + MEM[48571];
assign MEM[49187] = MEM[48511] + MEM[48577];
assign MEM[49188] = MEM[48512] + MEM[48580];
assign MEM[49189] = MEM[48513] + MEM[48565];
assign MEM[49190] = MEM[48514] + MEM[48574];
assign MEM[49191] = MEM[48515] + MEM[48581];
assign MEM[49192] = MEM[48516] + MEM[48576];
assign MEM[49193] = MEM[48518] + MEM[48572];
assign MEM[49194] = MEM[48522] + MEM[48592];
assign MEM[49195] = MEM[48523] + MEM[48600];
assign MEM[49196] = MEM[48526] + MEM[48610];
assign MEM[49197] = MEM[48527] + MEM[48570];
assign MEM[49198] = MEM[48529] + MEM[48594];
assign MEM[49199] = MEM[48530] + MEM[48606];
assign MEM[49200] = MEM[48531] + MEM[48584];
assign MEM[49201] = MEM[48536] + MEM[48604];
assign MEM[49202] = MEM[48538] + MEM[48579];
assign MEM[49203] = MEM[48539] + MEM[48624];
assign MEM[49204] = MEM[48544] + MEM[48573];
assign MEM[49205] = MEM[48545] + MEM[48598];
assign MEM[49206] = MEM[48548] + MEM[48619];
assign MEM[49207] = MEM[48549] + MEM[48637];
assign MEM[49208] = MEM[48550] + MEM[48607];
assign MEM[49209] = MEM[48552] + MEM[48608];
assign MEM[49210] = MEM[48553] + MEM[48620];
assign MEM[49211] = MEM[48554] + MEM[48597];
assign MEM[49212] = MEM[48558] + MEM[48609];
assign MEM[49213] = MEM[48559] + MEM[48616];
assign MEM[49214] = MEM[48561] + MEM[48617];
assign MEM[49215] = MEM[48562] + MEM[48638];
assign MEM[49216] = MEM[48563] + MEM[48629];
assign MEM[49217] = MEM[48566] + MEM[48649];
assign MEM[49218] = MEM[48567] + MEM[48633];
assign MEM[49219] = MEM[48568] + MEM[48623];
assign MEM[49220] = MEM[48582] + MEM[48642];
assign MEM[49221] = MEM[48583] + MEM[48639];
assign MEM[49222] = MEM[48585] + MEM[48666];
assign MEM[49223] = MEM[48586] + MEM[48654];
assign MEM[49224] = MEM[48587] + MEM[48645];
assign MEM[49225] = MEM[48588] + MEM[48660];
assign MEM[49226] = MEM[48589] + MEM[48653];
assign MEM[49227] = MEM[48590] + MEM[48656];
assign MEM[49228] = MEM[48591] + MEM[48644];
assign MEM[49229] = MEM[48593] + MEM[48640];
assign MEM[49230] = MEM[48595] + MEM[48661];
assign MEM[49231] = MEM[48596] + MEM[48655];
assign MEM[49232] = MEM[48599] + MEM[48692];
assign MEM[49233] = MEM[48601] + MEM[48659];
assign MEM[49234] = MEM[48602] + MEM[48643];
assign MEM[49235] = MEM[48603] + MEM[48658];
assign MEM[49236] = MEM[48605] + MEM[48647];
assign MEM[49237] = MEM[48611] + MEM[48682];
assign MEM[49238] = MEM[48612] + MEM[48672];
assign MEM[49239] = MEM[48613] + MEM[48678];
assign MEM[49240] = MEM[48614] + MEM[48696];
assign MEM[49241] = MEM[48615] + MEM[48681];
assign MEM[49242] = MEM[48618] + MEM[48676];
assign MEM[49243] = MEM[48621] + MEM[48686];
assign MEM[49244] = MEM[48622] + MEM[48703];
assign MEM[49245] = MEM[48625] + MEM[48683];
assign MEM[49246] = MEM[48626] + MEM[48699];
assign MEM[49247] = MEM[48627] + MEM[48685];
assign MEM[49248] = MEM[48628] + MEM[48711];
assign MEM[49249] = MEM[48630] + MEM[48679];
assign MEM[49250] = MEM[48631] + MEM[48700];
assign MEM[49251] = MEM[48632] + MEM[48695];
assign MEM[49252] = MEM[48634] + MEM[48690];
assign MEM[49253] = MEM[48635] + MEM[48704];
assign MEM[49254] = MEM[48636] + MEM[48688];
assign MEM[49255] = MEM[48641] + MEM[48691];
assign MEM[49256] = MEM[48646] + MEM[48725];
assign MEM[49257] = MEM[48648] + MEM[48734];
assign MEM[49258] = MEM[48650] + MEM[48702];
assign MEM[49259] = MEM[48651] + MEM[48706];
assign MEM[49260] = MEM[48652] + MEM[48737];
assign MEM[49261] = MEM[48657] + MEM[48729];
assign MEM[49262] = MEM[48662] + MEM[48736];
assign MEM[49263] = MEM[48663] + MEM[48731];
assign MEM[49264] = MEM[48664] + MEM[48709];
assign MEM[49265] = MEM[48665] + MEM[48744];
assign MEM[49266] = MEM[48667] + MEM[48712];
assign MEM[49267] = MEM[48668] + MEM[48738];
assign MEM[49268] = MEM[48669] + MEM[48762];
assign MEM[49269] = MEM[48670] + MEM[48727];
assign MEM[49270] = MEM[48671] + MEM[48716];
assign MEM[49271] = MEM[48673] + MEM[48720];
assign MEM[49272] = MEM[48674] + MEM[48735];
assign MEM[49273] = MEM[48675] + MEM[48717];
assign MEM[49274] = MEM[48677] + MEM[48764];
assign MEM[49275] = MEM[48680] + MEM[48754];
assign MEM[49276] = MEM[48684] + MEM[48740];
assign MEM[49277] = MEM[48687] + MEM[48767];
assign MEM[49278] = MEM[48689] + MEM[48749];
assign MEM[49279] = MEM[48693] + MEM[48745];
assign MEM[49280] = MEM[48694] + MEM[48760];
assign MEM[49281] = MEM[48697] + MEM[48765];
assign MEM[49282] = MEM[48698] + MEM[48774];
assign MEM[49283] = MEM[48701] + MEM[48757];
assign MEM[49284] = MEM[48705] + MEM[48759];
assign MEM[49285] = MEM[48707] + MEM[48756];
assign MEM[49286] = MEM[48708] + MEM[48752];
assign MEM[49287] = MEM[48710] + MEM[48769];
assign MEM[49288] = MEM[48713] + MEM[48781];
assign MEM[49289] = MEM[48714] + MEM[48793];
assign MEM[49290] = MEM[48715] + MEM[48777];
assign MEM[49291] = MEM[48718] + MEM[48779];
assign MEM[49292] = MEM[48719] + MEM[48802];
assign MEM[49293] = MEM[48721] + MEM[48796];
assign MEM[49294] = MEM[48722] + MEM[48780];
assign MEM[49295] = MEM[48723] + MEM[48795];
assign MEM[49296] = MEM[48724] + MEM[48817];
assign MEM[49297] = MEM[48726] + MEM[48798];
assign MEM[49298] = MEM[48728] + MEM[48790];
assign MEM[49299] = MEM[48730] + MEM[48801];
assign MEM[49300] = MEM[48732] + MEM[48800];
assign MEM[49301] = MEM[48733] + MEM[48792];
assign MEM[49302] = MEM[48739] + MEM[48782];
assign MEM[49303] = MEM[48741] + MEM[48814];
assign MEM[49304] = MEM[48742] + MEM[48799];
assign MEM[49305] = MEM[48743] + MEM[48804];
assign MEM[49306] = MEM[48746] + MEM[48812];
assign MEM[49307] = MEM[48747] + MEM[48807];
assign MEM[49308] = MEM[48748] + MEM[48813];
assign MEM[49309] = MEM[48750] + MEM[48787];
assign MEM[49310] = MEM[48751] + MEM[48806];
assign MEM[49311] = MEM[48753] + MEM[48857];
assign MEM[49312] = MEM[48755] + MEM[48794];
assign MEM[49313] = MEM[48758] + MEM[48815];
assign MEM[49314] = MEM[48761] + MEM[48820];
assign MEM[49315] = MEM[48763] + MEM[48830];
assign MEM[49316] = MEM[48766] + MEM[48847];
assign MEM[49317] = MEM[48768] + MEM[48826];
assign MEM[49318] = MEM[48770] + MEM[48832];
assign MEM[49319] = MEM[48771] + MEM[48833];
assign MEM[49320] = MEM[48772] + MEM[48848];
assign MEM[49321] = MEM[48773] + MEM[48824];
assign MEM[49322] = MEM[48775] + MEM[48851];
assign MEM[49323] = MEM[48776] + MEM[48839];
assign MEM[49324] = MEM[48778] + MEM[48837];
assign MEM[49325] = MEM[48783] + MEM[48842];
assign MEM[49326] = MEM[48784] + MEM[48856];
assign MEM[49327] = MEM[48785] + MEM[48828];
assign MEM[49328] = MEM[48786] + MEM[48855];
assign MEM[49329] = MEM[48788] + MEM[48861];
assign MEM[49330] = MEM[48789] + MEM[48868];
assign MEM[49331] = MEM[48791] + MEM[48850];
assign MEM[49332] = MEM[48797] + MEM[48831];
assign MEM[49333] = MEM[48803] + MEM[48863];
assign MEM[49334] = MEM[48805] + MEM[48864];
assign MEM[49335] = MEM[48808] + MEM[48870];
assign MEM[49336] = MEM[48809] + MEM[48871];
assign MEM[49337] = MEM[48810] + MEM[48872];
assign MEM[49338] = MEM[48811] + MEM[48877];
assign MEM[49339] = MEM[48816] + MEM[48878];
assign MEM[49340] = MEM[48818] + MEM[48898];
assign MEM[49341] = MEM[48819] + MEM[48879];
assign MEM[49342] = MEM[48821] + MEM[48885];
assign MEM[49343] = MEM[48822] + MEM[48852];
assign MEM[49344] = MEM[48823] + MEM[48889];
assign MEM[49345] = MEM[48825] + MEM[48887];
assign MEM[49346] = MEM[48827] + MEM[48902];
assign MEM[49347] = MEM[48829] + MEM[48892];
assign MEM[49348] = MEM[48834] + MEM[48912];
assign MEM[49349] = MEM[48835] + MEM[48895];
assign MEM[49350] = MEM[48836] + MEM[48900];
assign MEM[49351] = MEM[48838] + MEM[48881];
assign MEM[49352] = MEM[48840] + MEM[48928];
assign MEM[49353] = MEM[48841] + MEM[48914];
assign MEM[49354] = MEM[48843] + MEM[48911];
assign MEM[49355] = MEM[48844] + MEM[48929];
assign MEM[49356] = MEM[48845] + MEM[48901];
assign MEM[49357] = MEM[48846] + MEM[48917];
assign MEM[49358] = MEM[48849] + MEM[48893];
assign MEM[49359] = MEM[48853] + MEM[48915];
assign MEM[49360] = MEM[48854] + MEM[48924];
assign MEM[49361] = MEM[48858] + MEM[48904];
assign MEM[49362] = MEM[48859] + MEM[48907];
assign MEM[49363] = MEM[48860] + MEM[48923];
assign MEM[49364] = MEM[48862] + MEM[48930];
assign MEM[49365] = MEM[48865] + MEM[48908];
assign MEM[49366] = MEM[48866] + MEM[48935];
assign MEM[49367] = MEM[48867] + MEM[48936];
assign MEM[49368] = MEM[48869] + MEM[48938];
assign MEM[49369] = MEM[48873] + MEM[48942];
assign MEM[49370] = MEM[48874] + MEM[48894];
assign MEM[49371] = MEM[48875] + MEM[48913];
assign MEM[49372] = MEM[48876] + MEM[48934];
assign MEM[49373] = MEM[48880] + MEM[48945];
assign MEM[49374] = MEM[48882] + MEM[48952];
assign MEM[49375] = MEM[48883] + MEM[48969];
assign MEM[49376] = MEM[48884] + MEM[48933];
assign MEM[49377] = MEM[48886] + MEM[48954];
assign MEM[49378] = MEM[48888] + MEM[48932];
assign MEM[49379] = MEM[48890] + MEM[48956];
assign MEM[49380] = MEM[48891] + MEM[48949];
assign MEM[49381] = MEM[48896] + MEM[48950];
assign MEM[49382] = MEM[48897] + MEM[48966];
assign MEM[49383] = MEM[48899] + MEM[48992];
assign MEM[49384] = MEM[48903] + MEM[48980];
assign MEM[49385] = MEM[48905] + MEM[48974];
assign MEM[49386] = MEM[48906] + MEM[48970];
assign MEM[49387] = MEM[48909] + MEM[48964];
assign MEM[49388] = MEM[48910] + MEM[48957];
assign MEM[49389] = MEM[48916] + MEM[48986];
assign MEM[49390] = MEM[48918] + MEM[48968];
assign MEM[49391] = MEM[48919] + MEM[48979];
assign MEM[49392] = MEM[48920] + MEM[48987];
assign MEM[49393] = MEM[48921] + MEM[48982];
assign MEM[49394] = MEM[48922] + MEM[48996];
assign MEM[49395] = MEM[48925] + MEM[48976];
assign MEM[49396] = MEM[48926] + MEM[48990];
assign MEM[49397] = MEM[48927] + MEM[48984];
assign MEM[49398] = MEM[48931] + MEM[48997];
assign MEM[49399] = MEM[48937] + MEM[49034];
assign MEM[49400] = MEM[48939] + MEM[48998];
assign MEM[49401] = MEM[48940] + MEM[49011];
assign MEM[49402] = MEM[48941] + MEM[49028];
assign MEM[49403] = MEM[48943] + MEM[49015];
assign MEM[49404] = MEM[48944] + MEM[49005];
assign MEM[49405] = MEM[48946] + MEM[49030];
assign MEM[49406] = MEM[48947] + MEM[49031];
assign MEM[49407] = MEM[48948] + MEM[49016];
assign MEM[49408] = MEM[48951] + MEM[49007];
assign MEM[49409] = MEM[48953] + MEM[49000];
assign MEM[49410] = MEM[48955] + MEM[49017];
assign MEM[49411] = MEM[48958] + MEM[49020];
assign MEM[49412] = MEM[48959] + MEM[49035];
assign MEM[49413] = MEM[48960] + MEM[49018];
assign MEM[49414] = MEM[48961] + MEM[49008];
assign MEM[49415] = MEM[48962] + MEM[49027];
assign MEM[49416] = MEM[48963] + MEM[49013];
assign MEM[49417] = MEM[48965] + MEM[49024];
assign MEM[49418] = MEM[48967] + MEM[49019];
assign MEM[49419] = MEM[48971] + MEM[49042];
assign MEM[49420] = MEM[48972] + MEM[49047];
assign MEM[49421] = MEM[48973] + MEM[49040];
assign MEM[49422] = MEM[48975] + MEM[49025];
assign MEM[49423] = MEM[48977] + MEM[49022];
assign MEM[49424] = MEM[48978] + MEM[49029];
assign MEM[49425] = MEM[48981] + MEM[49033];
assign MEM[49426] = MEM[48983] + MEM[49036];
assign MEM[49427] = MEM[48985] + MEM[49032];
assign MEM[49428] = MEM[48988] + MEM[49051];
assign MEM[49429] = MEM[48989] + MEM[49041];
assign MEM[49430] = MEM[48991] + MEM[49068];
assign MEM[49431] = MEM[48993] + MEM[49067];
assign MEM[49432] = MEM[48994] + MEM[49048];
assign MEM[49433] = MEM[48995] + MEM[49058];
assign MEM[49434] = MEM[48999] + MEM[49094];
assign MEM[49435] = MEM[49001] + MEM[49050];
assign MEM[49436] = MEM[49002] + MEM[49066];
assign MEM[49437] = MEM[49003] + MEM[49056];
assign MEM[49438] = MEM[49004] + MEM[49071];
assign MEM[49439] = MEM[49006] + MEM[49069];
assign MEM[49440] = MEM[49009] + MEM[49057];
assign MEM[49441] = MEM[49010] + MEM[49095];
assign MEM[49442] = MEM[49012] + MEM[49070];
assign MEM[49443] = MEM[49014] + MEM[49083];
assign MEM[49444] = MEM[49021] + MEM[49076];
assign MEM[49445] = MEM[49023] + MEM[49096];
assign MEM[49446] = MEM[49026] + MEM[49072];
assign MEM[49447] = MEM[49037] + MEM[49079];
assign MEM[49448] = MEM[49038] + MEM[49089];
assign MEM[49449] = MEM[49039] + MEM[49080];
assign MEM[49450] = MEM[49043] + MEM[49123];
assign MEM[49451] = MEM[49044] + MEM[49112];
assign MEM[49452] = MEM[49045] + MEM[49110];
assign MEM[49453] = MEM[49046] + MEM[49117];
assign MEM[49454] = MEM[49049] + MEM[49119];
assign MEM[49455] = MEM[49052] + MEM[49132];
assign MEM[49456] = MEM[49053] + MEM[49134];
assign MEM[49457] = MEM[49054] + MEM[49121];
assign MEM[49458] = MEM[49055] + MEM[49125];
assign MEM[49459] = MEM[49059] + MEM[49147];
assign MEM[49460] = MEM[49060] + MEM[49127];
assign MEM[49461] = MEM[49061] + MEM[49131];
assign MEM[49462] = MEM[49062] + MEM[49122];
assign MEM[49463] = MEM[49063] + MEM[49116];
assign MEM[49464] = MEM[49064] + MEM[49113];
assign MEM[49465] = MEM[49065] + MEM[49139];
assign MEM[49466] = MEM[49073] + MEM[49166];
assign MEM[49467] = MEM[49074] + MEM[49168];
assign MEM[49468] = MEM[49075] + MEM[49124];
assign MEM[49469] = MEM[49077] + MEM[49173];
assign MEM[49470] = MEM[49078] + MEM[49136];
assign MEM[49471] = MEM[49081] + MEM[49145];
assign MEM[49472] = MEM[49082] + MEM[49141];
assign MEM[49473] = MEM[49084] + MEM[49154];
assign MEM[49474] = MEM[49085] + MEM[49153];
assign MEM[49475] = MEM[49086] + MEM[49144];
assign MEM[49476] = MEM[49087] + MEM[49151];
assign MEM[49477] = MEM[49088] + MEM[49155];
assign MEM[49478] = MEM[49090] + MEM[49146];
assign MEM[49479] = MEM[49091] + MEM[49152];
assign MEM[49480] = MEM[49092] + MEM[49160];
assign MEM[49481] = MEM[49093] + MEM[49158];
assign MEM[49482] = MEM[49097] + MEM[49161];
assign MEM[49483] = MEM[49098] + MEM[49157];
assign MEM[49484] = MEM[49099] + MEM[49150];
assign MEM[49485] = MEM[49100] + MEM[49181];
assign MEM[49486] = MEM[49101] + MEM[49163];
assign MEM[49487] = MEM[49102] + MEM[49156];
assign MEM[49488] = MEM[49103] + MEM[49165];
assign MEM[49489] = MEM[49104] + MEM[49164];
assign MEM[49490] = MEM[49105] + MEM[49172];
assign MEM[49491] = MEM[49106] + MEM[49167];
assign MEM[49492] = MEM[49107] + MEM[49176];
assign MEM[49493] = MEM[49108] + MEM[49170];
assign MEM[49494] = MEM[49109] + MEM[49180];
assign MEM[49495] = MEM[49111] + MEM[49169];
assign MEM[49496] = MEM[49114] + MEM[49179];
assign MEM[49497] = MEM[49115] + MEM[49175];
assign MEM[49498] = MEM[49118] + MEM[49177];
assign MEM[49499] = MEM[49120] + MEM[49183];
assign MEM[49500] = MEM[49126] + MEM[49182];
assign MEM[49501] = MEM[49128] + MEM[49193];
assign MEM[49502] = MEM[49129] + MEM[49178];
assign MEM[49503] = MEM[49130] + MEM[49205];
assign MEM[49504] = MEM[49133] + MEM[49196];
assign MEM[49505] = MEM[49135] + MEM[49189];
assign MEM[49506] = MEM[49137] + MEM[49186];
assign MEM[49507] = MEM[49138] + MEM[49187];
assign MEM[49508] = MEM[49140] + MEM[49191];
assign MEM[49509] = MEM[49142] + MEM[49199];
assign MEM[49510] = MEM[49143] + MEM[49204];
assign MEM[49511] = MEM[49148] + MEM[49202];
assign MEM[49512] = MEM[49149] + MEM[49197];
assign MEM[49513] = MEM[49159] + MEM[49212];
assign MEM[49514] = MEM[49162] + MEM[49242];
assign MEM[49515] = MEM[49171] + MEM[49246];
assign MEM[49516] = MEM[49174] + MEM[49221];
assign MEM[49517] = MEM[49184] + MEM[49259];
assign MEM[49518] = MEM[49185] + MEM[49253];
assign MEM[49519] = MEM[49188] + MEM[49263];
assign MEM[49520] = MEM[49190] + MEM[49271];
assign MEM[49521] = MEM[49192] + MEM[49244];
assign MEM[49522] = MEM[49194] + MEM[49257];
assign MEM[49523] = MEM[49195] + MEM[49272];
assign MEM[49524] = MEM[49198] + MEM[49261];
assign MEM[49525] = MEM[49200] + MEM[49258];
assign MEM[49526] = MEM[49201] + MEM[49260];
assign MEM[49527] = MEM[49203] + MEM[49280];
assign MEM[49528] = MEM[49206] + MEM[49276];
assign MEM[49529] = MEM[49207] + MEM[49278];
assign MEM[49530] = MEM[49208] + MEM[49270];
assign MEM[49531] = MEM[49209] + MEM[49269];
assign MEM[49532] = MEM[49210] + MEM[49286];
assign MEM[49533] = MEM[49211] + MEM[49266];
assign MEM[49534] = MEM[49213] + MEM[49268];
assign MEM[49535] = MEM[49214] + MEM[49262];
assign MEM[49536] = MEM[49215] + MEM[49285];
assign MEM[49537] = MEM[49216] + MEM[49279];
assign MEM[49538] = MEM[49217] + MEM[49290];
assign MEM[49539] = MEM[49218] + MEM[49282];
assign MEM[49540] = MEM[49219] + MEM[49274];
assign MEM[49541] = MEM[49220] + MEM[49287];
assign MEM[49542] = MEM[49222] + MEM[49300];
assign MEM[49543] = MEM[49223] + MEM[49295];
assign MEM[49544] = MEM[49224] + MEM[49284];
assign MEM[49545] = MEM[49225] + MEM[49292];
assign MEM[49546] = MEM[49226] + MEM[49293];
assign MEM[49547] = MEM[49227] + MEM[49288];
assign MEM[49548] = MEM[49228] + MEM[49281];
assign MEM[49549] = MEM[49229] + MEM[49283];
assign MEM[49550] = MEM[49230] + MEM[49298];
assign MEM[49551] = MEM[49231] + MEM[49296];
assign MEM[49552] = MEM[49232] + MEM[49291];
assign MEM[49553] = MEM[49233] + MEM[49307];
assign MEM[49554] = MEM[49234] + MEM[49304];
assign MEM[49555] = MEM[49235] + MEM[49299];
assign MEM[49556] = MEM[49236] + MEM[49305];
assign MEM[49557] = MEM[49237] + MEM[49302];
assign MEM[49558] = MEM[49238] + MEM[49297];
assign MEM[49559] = MEM[49239] + MEM[49312];
assign MEM[49560] = MEM[49240] + MEM[49309];
assign MEM[49561] = MEM[49241] + MEM[49294];
assign MEM[49562] = MEM[49243] + MEM[49310];
assign MEM[49563] = MEM[49245] + MEM[49314];
assign MEM[49564] = MEM[49247] + MEM[49301];
assign MEM[49565] = MEM[49248] + MEM[49317];
assign MEM[49566] = MEM[49249] + MEM[49308];
assign MEM[49567] = MEM[49250] + MEM[49315];
assign MEM[49568] = MEM[49251] + MEM[49306];
assign MEM[49569] = MEM[49252] + MEM[49318];
assign MEM[49570] = MEM[49254] + MEM[49303];
assign MEM[49571] = MEM[49255] + MEM[49319];
assign MEM[49572] = MEM[49256] + MEM[49331];
assign MEM[49573] = MEM[49264] + MEM[49311];
assign MEM[49574] = MEM[49265] + MEM[49316];
assign MEM[49575] = MEM[49267] + MEM[49336];
assign MEM[49576] = MEM[49273] + MEM[49326];
assign MEM[49577] = MEM[49275] + MEM[49343];
assign MEM[49578] = MEM[49277] + MEM[49349];
assign MEM[49579] = MEM[49289] + MEM[49370];
assign MEM[49580] = MEM[49313] + MEM[49373];
assign MEM[49581] = MEM[49320] + MEM[49402];
assign MEM[49582] = MEM[49321] + MEM[49375];
assign MEM[49583] = MEM[49322] + MEM[49398];
assign MEM[49584] = MEM[49323] + MEM[49397];
assign MEM[49585] = MEM[49324] + MEM[49382];
assign MEM[49586] = MEM[49325] + MEM[49387];
assign MEM[49587] = MEM[49327] + MEM[49383];
assign MEM[49588] = MEM[49328] + MEM[49392];
assign MEM[49589] = MEM[49329] + MEM[49391];
assign MEM[49590] = MEM[49330] + MEM[49401];
assign MEM[49591] = MEM[49332] + MEM[49395];
assign MEM[49592] = MEM[49333] + MEM[49396];
assign MEM[49593] = MEM[49334] + MEM[49389];
assign MEM[49594] = MEM[49335] + MEM[49400];
assign MEM[49595] = MEM[49337] + MEM[49403];
assign MEM[49596] = MEM[49338] + MEM[49404];
assign MEM[49597] = MEM[49339] + MEM[49409];
assign MEM[49598] = MEM[49340] + MEM[49418];
assign MEM[49599] = MEM[49341] + MEM[49408];
assign MEM[49600] = MEM[49342] + MEM[49416];
assign MEM[49601] = MEM[49344] + MEM[49413];
assign MEM[49602] = MEM[49345] + MEM[49399];
assign MEM[49603] = MEM[49346] + MEM[49427];
assign MEM[49604] = MEM[49347] + MEM[49407];
assign MEM[49605] = MEM[49348] + MEM[49421];
assign MEM[49606] = MEM[49350] + MEM[49405];
assign MEM[49607] = MEM[49351] + MEM[49415];
assign MEM[49608] = MEM[49352] + MEM[49428];
assign MEM[49609] = MEM[49353] + MEM[49425];
assign MEM[49610] = MEM[49354] + MEM[49406];
assign MEM[49611] = MEM[49355] + MEM[49432];
assign MEM[49612] = MEM[49356] + MEM[49422];
assign MEM[49613] = MEM[49357] + MEM[49420];
assign MEM[49614] = MEM[49358] + MEM[49412];
assign MEM[49615] = MEM[49359] + MEM[49423];
assign MEM[49616] = MEM[49360] + MEM[49438];
assign MEM[49617] = MEM[49361] + MEM[49411];
assign MEM[49618] = MEM[49362] + MEM[49426];
assign MEM[49619] = MEM[49363] + MEM[49424];
assign MEM[49620] = MEM[49364] + MEM[49439];
assign MEM[49621] = MEM[49365] + MEM[49417];
assign MEM[49622] = MEM[49366] + MEM[49430];
assign MEM[49623] = MEM[49367] + MEM[49433];
assign MEM[49624] = MEM[49368] + MEM[49436];
assign MEM[49625] = MEM[49369] + MEM[49429];
assign MEM[49626] = MEM[49371] + MEM[49419];
assign MEM[49627] = MEM[49372] + MEM[49434];
assign MEM[49628] = MEM[49374] + MEM[49443];
assign MEM[49629] = MEM[49376] + MEM[49441];
assign MEM[49630] = MEM[49377] + MEM[49440];
assign MEM[49631] = MEM[49378] + MEM[49431];
assign MEM[49632] = MEM[49379] + MEM[49437];
assign MEM[49633] = MEM[49380] + MEM[49442];
assign MEM[49634] = MEM[49381] + MEM[49435];
assign MEM[49635] = MEM[49384] + MEM[49449];
assign MEM[49636] = MEM[49385] + MEM[49448];
assign MEM[49637] = MEM[49386] + MEM[49444];
assign MEM[49638] = MEM[49388] + MEM[49447];
assign MEM[49639] = MEM[49390] + MEM[49445];
assign MEM[49640] = MEM[49393] + MEM[49446];
assign MEM[49641] = MEM[49394] + MEM[49469];
assign MEM[49642] = MEM[49410] + MEM[49464];
assign MEM[49643] = MEM[49414] + MEM[49463];
assign MEM[49644] = MEM[49450] + MEM[49523];
assign MEM[49645] = MEM[49451] + MEM[49522];
assign MEM[49646] = MEM[49452] + MEM[49515];
assign MEM[49647] = MEM[49453] + MEM[49519];
assign MEM[49648] = MEM[49454] + MEM[49521];
assign MEM[49649] = MEM[49455] + MEM[49520];
assign MEM[49650] = MEM[49456] + MEM[49531];
assign MEM[49651] = MEM[49457] + MEM[49517];
assign MEM[49652] = MEM[49458] + MEM[49525];
assign MEM[49653] = MEM[49459] + MEM[49533];
assign MEM[49654] = MEM[49460] + MEM[49518];
assign MEM[49655] = MEM[49461] + MEM[49537];
assign MEM[49656] = MEM[49462] + MEM[49524];
assign MEM[49657] = MEM[49465] + MEM[49532];
assign MEM[49658] = MEM[49466] + MEM[49535];
assign MEM[49659] = MEM[49467] + MEM[49544];
assign MEM[49660] = MEM[49468] + MEM[49528];
assign MEM[49661] = MEM[49470] + MEM[49526];
assign MEM[49662] = MEM[49471] + MEM[49536];
assign MEM[49663] = MEM[49472] + MEM[49534];
assign MEM[49664] = MEM[49473] + MEM[49545];
assign MEM[49665] = MEM[49474] + MEM[49538];
assign MEM[49666] = MEM[49475] + MEM[49530];
assign MEM[49667] = MEM[49476] + MEM[49527];
assign MEM[49668] = MEM[49477] + MEM[49559];
assign MEM[49669] = MEM[49478] + MEM[49539];
assign MEM[49670] = MEM[49479] + MEM[49547];
assign MEM[49671] = MEM[49480] + MEM[49546];
assign MEM[49672] = MEM[49481] + MEM[49529];
assign MEM[49673] = MEM[49482] + MEM[49549];
assign MEM[49674] = MEM[49483] + MEM[49551];
assign MEM[49675] = MEM[49484] + MEM[49541];
assign MEM[49676] = MEM[49485] + MEM[49560];
assign MEM[49677] = MEM[49486] + MEM[49542];
assign MEM[49678] = MEM[49487] + MEM[49543];
assign MEM[49679] = MEM[49488] + MEM[49556];
assign MEM[49680] = MEM[49489] + MEM[49548];
assign MEM[49681] = MEM[49490] + MEM[49554];
assign MEM[49682] = MEM[49491] + MEM[49550];
assign MEM[49683] = MEM[49492] + MEM[49564];
assign MEM[49684] = MEM[49493] + MEM[49567];
assign MEM[49685] = MEM[49494] + MEM[49552];
assign MEM[49686] = MEM[49495] + MEM[49540];
assign MEM[49687] = MEM[49496] + MEM[49553];
assign MEM[49688] = MEM[49497] + MEM[49562];
assign MEM[49689] = MEM[49498] + MEM[49565];
assign MEM[49690] = MEM[49499] + MEM[49555];
assign MEM[49691] = MEM[49500] + MEM[49557];
assign MEM[49692] = MEM[49501] + MEM[49568];
assign MEM[49693] = MEM[49502] + MEM[49561];
assign MEM[49694] = MEM[49503] + MEM[49573];
assign MEM[49695] = MEM[49504] + MEM[49575];
assign MEM[49696] = MEM[49505] + MEM[49570];
assign MEM[49697] = MEM[49506] + MEM[49558];
assign MEM[49698] = MEM[49507] + MEM[49563];
assign MEM[49699] = MEM[49508] + MEM[49572];
assign MEM[49700] = MEM[49509] + MEM[49574];
assign MEM[49701] = MEM[49510] + MEM[49566];
assign MEM[49702] = MEM[49511] + MEM[49571];
assign MEM[49703] = MEM[49512] + MEM[49569];
assign MEM[49704] = MEM[49513] + MEM[49576];
assign MEM[49705] = MEM[49514] + MEM[49579];
assign MEM[49706] = MEM[49516] + MEM[49578];
assign MEM[49707] = MEM[49577] + MEM[49641];
assign MEM[49708] = MEM[49580] + MEM[49648];
assign MEM[49709] = MEM[49581] + MEM[49666];
assign MEM[49710] = MEM[49582] + MEM[49646];
assign MEM[49711] = MEM[49583] + MEM[49654];
assign MEM[49712] = MEM[49584] + MEM[49651];
assign MEM[49713] = MEM[49585] + MEM[49647];
assign MEM[49714] = MEM[49586] + MEM[49649];
assign MEM[49715] = MEM[49587] + MEM[49652];
assign MEM[49716] = MEM[49588] + MEM[49656];
assign MEM[49717] = MEM[49589] + MEM[49644];
assign MEM[49718] = MEM[49590] + MEM[49660];
assign MEM[49719] = MEM[49591] + MEM[49645];
assign MEM[49720] = MEM[49592] + MEM[49661];
assign MEM[49721] = MEM[49593] + MEM[49650];
assign MEM[49722] = MEM[49594] + MEM[49653];
assign MEM[49723] = MEM[49595] + MEM[49658];
assign MEM[49724] = MEM[49596] + MEM[49655];
assign MEM[49725] = MEM[49597] + MEM[49657];
assign MEM[49726] = MEM[49598] + MEM[49659];
assign MEM[49727] = MEM[49599] + MEM[49663];
assign MEM[49728] = MEM[49600] + MEM[49672];
assign MEM[49729] = MEM[49601] + MEM[49667];
assign MEM[49730] = MEM[49602] + MEM[49686];
assign MEM[49731] = MEM[49603] + MEM[49673];
assign MEM[49732] = MEM[49604] + MEM[49665];
assign MEM[49733] = MEM[49605] + MEM[49685];
assign MEM[49734] = MEM[49606] + MEM[49680];
assign MEM[49735] = MEM[49607] + MEM[49662];
assign MEM[49736] = MEM[49608] + MEM[49682];
assign MEM[49737] = MEM[49609] + MEM[49671];
assign MEM[49738] = MEM[49610] + MEM[49681];
assign MEM[49739] = MEM[49611] + MEM[49678];
assign MEM[49740] = MEM[49612] + MEM[49664];
assign MEM[49741] = MEM[49613] + MEM[49679];
assign MEM[49742] = MEM[49614] + MEM[49669];
assign MEM[49743] = MEM[49615] + MEM[49670];
assign MEM[49744] = MEM[49616] + MEM[49693];
assign MEM[49745] = MEM[49617] + MEM[49675];
assign MEM[49746] = MEM[49618] + MEM[49668];
assign MEM[49747] = MEM[49619] + MEM[49677];
assign MEM[49748] = MEM[49620] + MEM[49687];
assign MEM[49749] = MEM[49621] + MEM[49674];
assign MEM[49750] = MEM[49622] + MEM[49691];
assign MEM[49751] = MEM[49623] + MEM[49690];
assign MEM[49752] = MEM[49624] + MEM[49697];
assign MEM[49753] = MEM[49625] + MEM[49676];
assign MEM[49754] = MEM[49626] + MEM[49688];
assign MEM[49755] = MEM[49627] + MEM[49701];
assign MEM[49756] = MEM[49628] + MEM[49696];
assign MEM[49757] = MEM[49629] + MEM[49703];
assign MEM[49758] = MEM[49630] + MEM[49683];
assign MEM[49759] = MEM[49631] + MEM[49698];
assign MEM[49760] = MEM[49632] + MEM[49689];
assign MEM[49761] = MEM[49633] + MEM[49692];
assign MEM[49762] = MEM[49634] + MEM[49684];
assign MEM[49763] = MEM[49635] + MEM[49699];
assign MEM[49764] = MEM[49636] + MEM[49700];
assign MEM[49765] = MEM[49637] + MEM[49694];
assign MEM[49766] = MEM[49638] + MEM[49702];
assign MEM[49767] = MEM[49639] + MEM[49704];
assign MEM[49768] = MEM[49640] + MEM[49695];
assign MEM[49769] = MEM[49642] + MEM[49705];
assign MEM[49770] = MEM[49643] + MEM[49706];
assign output_vector[0] = MEM[49710];
assign output_vector[1] = MEM[49723];
assign output_vector[2] = MEM[49713];
assign output_vector[3] = MEM[49758];
assign output_vector[4] = MEM[49748];
assign output_vector[5] = MEM[49725];
assign output_vector[6] = MEM[49737];
assign output_vector[7] = MEM[49714];
assign output_vector[8] = MEM[49759];
assign output_vector[9] = MEM[49761];
assign output_vector[10] = MEM[49764];
assign output_vector[11] = MEM[49766];
assign output_vector[12] = MEM[49709];
assign output_vector[13] = MEM[49756];
assign output_vector[14] = MEM[49732];
assign output_vector[15] = MEM[49762];
assign output_vector[16] = MEM[49754];
assign output_vector[17] = MEM[49717];
assign output_vector[18] = MEM[49738];
assign output_vector[19] = MEM[49752];
assign output_vector[20] = MEM[49745];
assign output_vector[21] = MEM[49746];
assign output_vector[22] = MEM[49755];
assign output_vector[23] = MEM[49731];
assign output_vector[24] = MEM[49739];
assign output_vector[25] = MEM[49749];
assign output_vector[26] = MEM[49721];
assign output_vector[27] = MEM[49751];
assign output_vector[28] = MEM[49707];
assign output_vector[29] = MEM[49722];
assign output_vector[30] = MEM[49743];
assign output_vector[31] = MEM[49765];
assign output_vector[32] = MEM[49711];
assign output_vector[33] = MEM[49720];
assign output_vector[34] = MEM[49730];
assign output_vector[35] = MEM[49763];
assign output_vector[36] = MEM[49767];
assign output_vector[37] = MEM[49742];
assign output_vector[38] = MEM[49741];
assign output_vector[39] = MEM[49747];
assign output_vector[40] = MEM[49729];
assign output_vector[41] = MEM[49734];
assign output_vector[42] = MEM[49753];
assign output_vector[43] = MEM[49736];
assign output_vector[44] = MEM[49757];
assign output_vector[45] = MEM[49708];
assign output_vector[46] = MEM[49728];
assign output_vector[47] = MEM[49726];
assign output_vector[48] = MEM[49719];
assign output_vector[49] = MEM[49712];
assign output_vector[50] = MEM[49727];
assign output_vector[51] = MEM[49715];
assign output_vector[52] = MEM[49770];
assign output_vector[53] = MEM[49724];
assign output_vector[54] = MEM[49744];
assign output_vector[55] = MEM[49740];
assign output_vector[56] = MEM[49750];
assign output_vector[57] = MEM[49735];
assign output_vector[58] = MEM[49769];
assign output_vector[59] = MEM[49733];
assign output_vector[60] = MEM[49768];
assign output_vector[61] = MEM[49760];
assign output_vector[62] = MEM[49716];
assign output_vector[63] = MEM[49718];

endmodule
